* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : bias                                         *
* Netlisted  : Mon Aug 26 08:37:01 2024                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(ne3) nem ndiff(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 1 MP(pe3) pem pdiff(D) p1trm(G) pdiff(S) nwtrm(B)
*.DEVTMPLT 2 NE3I_6() nemi_6 ndiff(D) p1trm(G) ndiff(S) pwitrm(B) dnwtrm(NW) bulk(SB)
*.DEVTMPLT 3 MOSVC3() mosvcm p1trm(G) nwtrm(NW) bulk(SB)
*.DEVTMPLT 4 Q(qpvc3) qpvmc bulk(C) nwtrm(B) pdiff(E)
*.DEVTMPLT 5 D(p_dnw) p_dnw bulk(POS) nwtrm(NEG)
*.DEVTMPLT 6 D(p_ddnw) p_ddnw bulk(POS) dnwtrm(NEG)
*.DEVTMPLT 7 D(p_dipdnwmv) p_dipwmv pwitrm(POS) dnwtrm(NEG)
*.DEVTMPLT 8 D(p_dnw3) p_dnwm bulk(POS) nwtrm(NEG)
*.DEVTMPLT 9 R(rpp1k1_3) rpp1k1_s p1trm(POS) p1trm(NEG) bulk(SUB)
*.DEVTMPLT 10 R(rpp1k1_3) rpp1k1_n p1trm(POS) p1trm(NEG) nwtrm(SUB)
*.DEVTMPLT 11 C(cmm5t) cmim capm(POS) m4trm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_724654214590                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_724654214590 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_724654214590

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_724654214593                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_724654214593 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_724654214593

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724654214594                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724654214594 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724654214594

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_724654214595                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_724654214595 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_724654214595

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724654214597                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724654214597 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724654214597

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724654214598                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724654214598 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724654214598

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724654214599                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724654214599 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724654214599

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246542145910                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246542145910 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246542145910

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246542145911                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246542145911 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246542145911

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246542145912                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246542145912 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246542145912

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246542145913                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246542145913 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246542145913

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246542145914                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246542145914 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246542145914

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246542145915                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246542145915 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246542145915

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246542145916                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246542145916 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246542145916

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246542145917                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246542145917 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246542145917

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246542145918                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246542145918 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246542145918

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246542145919                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246542145919 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246542145919

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246542145920                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246542145920 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246542145920

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246542145921                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246542145921 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246542145921

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246542145922                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246542145922 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246542145922

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246542145923                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246542145923 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246542145923

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246542145924                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246542145924 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246542145924

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_7246542145925                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_7246542145925 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_7246542145925

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246542145926                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246542145926 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246542145926

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246542145927                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246542145927 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246542145927

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246542145928                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246542145928 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246542145928

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246542145936                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246542145936 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246542145936

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246542145937                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246542145937 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246542145937

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246542145940                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246542145940 1 2
** N=2 EP=2 FDC=0
.ends VIA1_C_CDNS_7246542145940

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724654214590                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724654214590 1 2 3 4 5
** N=5 EP=5 FDC=11
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=1
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=1
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=1
M4 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=6160 $Y=0 $dt=1
M5 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7700 $Y=0 $dt=1
M6 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=9240 $Y=0 $dt=1
M7 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10780 $Y=0 $dt=1
M8 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12320 $Y=0 $dt=1
M9 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=13860 $Y=0 $dt=1
D10 5 4 p_dnw3 AREA=2.15633e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=8
.ends pe3_CDNS_724654214590

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724654214591                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724654214591 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
.ends ne3_CDNS_724654214591

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724654214592                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724654214592 1 2 3 4 5
** N=5 EP=5 FDC=13
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=1
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=1
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=1
M4 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=6160 $Y=0 $dt=1
M5 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7700 $Y=0 $dt=1
M6 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=9240 $Y=0 $dt=1
M7 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10780 $Y=0 $dt=1
M8 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12320 $Y=0 $dt=1
M9 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=13860 $Y=0 $dt=1
M10 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=15400 $Y=0 $dt=1
M11 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=16940 $Y=0 $dt=1
D12 5 4 p_dnw3 AREA=2.52778e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=8
.ends pe3_CDNS_724654214592

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724654214593                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724654214593 1 2 3 4
** N=4 EP=4 FDC=3
M0 2 2 1 3 pe3 L=2e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 2 3 pe3 L=2e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=2540 $Y=0 $dt=1
D2 4 3 p_dnw3 AREA=9.11736e-11 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=8
.ends pe3_CDNS_724654214593

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_724654214594                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_724654214594 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.0005141 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=9
.ends rpp1k1_3_CDNS_724654214594

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724654214595                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724654214595 1 2 3 4
** N=4 EP=4 FDC=8
M0 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
M1 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=2540 $Y=0 $dt=0
M2 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=5080 $Y=0 $dt=0
M3 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7620 $Y=0 $dt=0
M4 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10160 $Y=0 $dt=0
M5 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12700 $Y=0 $dt=0
M6 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=15240 $Y=0 $dt=0
M7 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=17780 $Y=0 $dt=0
.ends ne3_CDNS_724654214595

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724654214599                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724654214599 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
M0 3 2 1 1 pe3 L=2e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_724654214599

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246542145910                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246542145910 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
M0 3 2 1 1 pe3 L=1e-05 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_7246542145910

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3i_6_CDNS_724654214598                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3i_6_CDNS_724654214598 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=1
X0 1 2 3 1 4 5 NE3I_6 w=1e-05 l=2e-06 as=4.8e-12 ad=4.8e-12 ps=2.096e-05 pd=2.096e-05 $X=0 $Y=0 $dt=2
.ends ne3i_6_CDNS_724654214598

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A3                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A3 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=2
X0 1 4 5 6 7 ne3i_6_CDNS_724654214598 $T=4060 14570 1 0 $X=0 $Y=0
X1 1 2 3 6 7 ne3i_6_CDNS_724654214598 $T=7460 14570 1 0 $X=3400 $Y=0
.ends MASCO__A3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A4                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A4 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=2
X0 1 4 5 6 7 ne3i_6_CDNS_724654214598 $T=4060 4450 0 0 $X=0 $Y=0
X1 1 2 3 6 7 ne3i_6_CDNS_724654214598 $T=7460 4450 0 0 $X=3400 $Y=0
.ends MASCO__A4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__B5                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__B5 1 2 3 4 5 6 7 8 9 10
+ 11
*.DEVICECLIMB
** N=11 EP=11 FDC=4
X0 1 10 6 5 3 2 11 MASCO__A3 $T=0 14680 0 0 $X=0 $Y=14680
X1 1 8 7 9 4 2 11 MASCO__A4 $T=0 0 0 0 $X=0 $Y=0
.ends MASCO__B5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ref_bias                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ref_bias 1 2 3 4 5 6 7
** N=18 EP=7 FDC=187
X0 8 VIA2_C_CDNS_724654214590 $T=152805 186425 0 0 $X=152055 $Y=185675
X1 5 VIA2_C_CDNS_724654214590 $T=187300 141530 0 0 $X=186550 $Y=140780
X2 9 VIA2_C_CDNS_724654214593 $T=13870 9200 0 0 $X=13160 $Y=8800
X3 9 VIA2_C_CDNS_724654214593 $T=13870 25290 0 0 $X=13160 $Y=24890
X4 8 VIA2_C_CDNS_724654214593 $T=64530 11760 0 0 $X=63820 $Y=11360
X5 8 VIA2_C_CDNS_724654214593 $T=64530 27850 0 0 $X=63820 $Y=27450
X6 10 VIA2_C_CDNS_724654214593 $T=66310 10480 0 0 $X=65600 $Y=10080
X7 10 VIA2_C_CDNS_724654214593 $T=66310 26570 0 0 $X=65600 $Y=26170
X8 1 VIA1_C_CDNS_724654214594 $T=17710 13040 0 0 $X=17570 $Y=12590
X9 1 VIA1_C_CDNS_724654214594 $T=17710 29130 0 0 $X=17570 $Y=28680
X10 1 VIA1_C_CDNS_724654214594 $T=20480 29130 0 0 $X=20340 $Y=28680
X11 1 VIA1_C_CDNS_724654214594 $T=20480 42300 0 0 $X=20340 $Y=41850
X12 1 VIA1_C_CDNS_724654214594 $T=23250 13040 0 0 $X=23110 $Y=12590
X13 1 VIA1_C_CDNS_724654214594 $T=23250 29130 0 0 $X=23110 $Y=28680
X14 1 VIA1_C_CDNS_724654214594 $T=23950 13040 0 0 $X=23810 $Y=12590
X15 1 VIA1_C_CDNS_724654214594 $T=23950 29130 0 0 $X=23810 $Y=28680
X16 9 VIA1_C_CDNS_724654214594 $T=26720 25290 0 0 $X=26580 $Y=24840
X17 10 VIA1_C_CDNS_724654214594 $T=29490 10480 0 0 $X=29350 $Y=10030
X18 9 VIA1_C_CDNS_724654214594 $T=29490 25290 0 0 $X=29350 $Y=24840
X19 1 VIA1_C_CDNS_724654214594 $T=30190 13040 0 0 $X=30050 $Y=12590
X20 1 VIA1_C_CDNS_724654214594 $T=30190 29130 0 0 $X=30050 $Y=28680
X21 9 VIA1_C_CDNS_724654214594 $T=32960 25290 0 0 $X=32820 $Y=24840
X22 9 VIA1_C_CDNS_724654214594 $T=35730 9200 0 0 $X=35590 $Y=8750
X23 10 VIA1_C_CDNS_724654214594 $T=35730 26570 0 0 $X=35590 $Y=26120
X24 1 VIA1_C_CDNS_724654214594 $T=36430 13040 0 0 $X=36290 $Y=12590
X25 1 VIA1_C_CDNS_724654214594 $T=36430 29130 0 0 $X=36290 $Y=28680
X26 9 VIA1_C_CDNS_724654214594 $T=39200 25290 0 0 $X=39060 $Y=24840
X27 8 VIA1_C_CDNS_724654214594 $T=41970 11760 0 0 $X=41830 $Y=11310
X28 9 VIA1_C_CDNS_724654214594 $T=41970 25290 0 0 $X=41830 $Y=24840
X29 1 VIA1_C_CDNS_724654214594 $T=42670 13040 0 0 $X=42530 $Y=12590
X30 1 VIA1_C_CDNS_724654214594 $T=42670 29130 0 0 $X=42530 $Y=28680
X31 9 VIA1_C_CDNS_724654214594 $T=45440 25290 0 0 $X=45300 $Y=24840
X32 9 VIA1_C_CDNS_724654214594 $T=48210 9200 0 0 $X=48070 $Y=8750
X33 10 VIA1_C_CDNS_724654214594 $T=48210 26570 0 0 $X=48070 $Y=26120
X34 1 VIA1_C_CDNS_724654214594 $T=48910 13040 0 0 $X=48770 $Y=12590
X35 1 VIA1_C_CDNS_724654214594 $T=48910 29130 0 0 $X=48770 $Y=28680
X36 9 VIA1_C_CDNS_724654214594 $T=51680 25290 0 0 $X=51540 $Y=24840
X37 1 VIA1_C_CDNS_724654214594 $T=51680 42300 0 0 $X=51540 $Y=41850
X38 10 VIA1_C_CDNS_724654214594 $T=54450 10480 0 0 $X=54310 $Y=10030
X39 1 VIA1_C_CDNS_724654214594 $T=54450 29130 0 0 $X=54310 $Y=28680
X40 1 VIA1_C_CDNS_724654214594 $T=55150 13040 0 0 $X=55010 $Y=12590
X41 1 VIA1_C_CDNS_724654214594 $T=55150 29130 0 0 $X=55010 $Y=28680
X42 1 VIA1_C_CDNS_724654214594 $T=57920 29130 0 0 $X=57780 $Y=28680
X43 1 VIA1_C_CDNS_724654214594 $T=57920 42300 0 0 $X=57780 $Y=41850
X44 1 VIA1_C_CDNS_724654214594 $T=60690 13040 0 0 $X=60550 $Y=12590
X45 1 VIA1_C_CDNS_724654214594 $T=60690 29130 0 0 $X=60550 $Y=28680
X46 1 VIA2_C_CDNS_724654214595 $T=15900 13040 0 0 $X=14930 $Y=12640
X47 1 VIA2_C_CDNS_724654214595 $T=15900 29130 0 0 $X=14930 $Y=28730
X48 1 VIA2_C_CDNS_724654214595 $T=15900 42300 0 0 $X=14930 $Y=41900
X49 1 VIA2_C_CDNS_724654214595 $T=62500 13040 0 0 $X=61530 $Y=12640
X50 1 VIA2_C_CDNS_724654214595 $T=62500 29130 0 0 $X=61530 $Y=28730
X51 1 VIA2_C_CDNS_724654214595 $T=62500 42300 0 0 $X=61530 $Y=41900
X52 9 VIA1_C_CDNS_724654214597 $T=26720 41270 0 0 $X=26580 $Y=41080
X53 9 VIA1_C_CDNS_724654214597 $T=32960 41270 0 0 $X=32820 $Y=41080
X54 9 VIA1_C_CDNS_724654214597 $T=39200 41270 0 0 $X=39060 $Y=41080
X55 9 VIA1_C_CDNS_724654214597 $T=45440 41270 0 0 $X=45300 $Y=41080
X56 9 VIA1_C_CDNS_724654214598 $T=17275 53125 0 0 $X=16875 $Y=52415
X57 3 VIA1_C_CDNS_724654214598 $T=19815 51345 0 0 $X=19415 $Y=50635
X58 9 VIA1_C_CDNS_724654214598 $T=22355 53125 0 0 $X=21955 $Y=52415
X59 3 VIA1_C_CDNS_724654214598 $T=24895 51345 0 0 $X=24495 $Y=50635
X60 9 VIA1_C_CDNS_724654214598 $T=27435 53125 0 0 $X=27035 $Y=52415
X61 3 VIA1_C_CDNS_724654214598 $T=29975 51345 0 0 $X=29575 $Y=50635
X62 9 VIA1_C_CDNS_724654214598 $T=32515 53125 0 0 $X=32115 $Y=52415
X63 3 VIA1_C_CDNS_724654214598 $T=35055 51345 0 0 $X=34655 $Y=50635
X64 9 VIA1_C_CDNS_724654214598 $T=37595 53125 0 0 $X=37195 $Y=52415
X65 10 VIA1_C_CDNS_724654214598 $T=42210 52905 0 0 $X=41810 $Y=52195
X66 11 VIA1_C_CDNS_724654214598 $T=44750 51125 0 0 $X=44350 $Y=50415
X67 10 VIA1_C_CDNS_724654214598 $T=47290 52905 0 0 $X=46890 $Y=52195
X68 11 VIA1_C_CDNS_724654214598 $T=49830 51125 0 0 $X=49430 $Y=50415
X69 10 VIA1_C_CDNS_724654214598 $T=52370 52905 0 0 $X=51970 $Y=52195
X70 11 VIA1_C_CDNS_724654214598 $T=54910 51125 0 0 $X=54510 $Y=50415
X71 10 VIA1_C_CDNS_724654214598 $T=57450 52905 0 0 $X=57050 $Y=52195
X72 11 VIA1_C_CDNS_724654214598 $T=59990 51125 0 0 $X=59590 $Y=50415
X73 10 VIA1_C_CDNS_724654214598 $T=62530 52905 0 0 $X=62130 $Y=52195
X74 2 VIA1_C_CDNS_724654214598 $T=137790 186425 0 0 $X=137390 $Y=185715
X75 12 VIA1_C_CDNS_724654214598 $T=140330 188205 0 0 $X=139930 $Y=187495
X76 2 VIA1_C_CDNS_724654214598 $T=142870 186425 0 0 $X=142470 $Y=185715
X77 12 VIA1_C_CDNS_724654214598 $T=147350 188205 0 0 $X=146950 $Y=187495
X78 8 VIA1_C_CDNS_724654214598 $T=149890 186425 0 0 $X=149490 $Y=185715
X79 12 VIA1_C_CDNS_724654214598 $T=152430 188205 0 0 $X=152030 $Y=187495
X80 13 VIA1_C_CDNS_724654214598 $T=162070 148400 0 0 $X=161670 $Y=147690
X81 4 VIA1_C_CDNS_724654214598 $T=163610 146620 0 0 $X=163210 $Y=145910
X82 13 VIA1_C_CDNS_724654214598 $T=165150 148400 0 0 $X=164750 $Y=147690
X83 2 VIA1_C_CDNS_724654214598 $T=165405 173875 0 0 $X=165005 $Y=173165
X84 2 VIA1_C_CDNS_724654214598 $T=165405 193895 0 0 $X=165005 $Y=193185
X85 2 VIA1_C_CDNS_724654214598 $T=166675 193895 0 0 $X=166275 $Y=193185
X86 2 VIA1_C_CDNS_724654214598 $T=166675 208575 0 0 $X=166275 $Y=207865
X87 4 VIA1_C_CDNS_724654214598 $T=166690 146620 0 0 $X=166290 $Y=145910
X88 2 VIA1_C_CDNS_724654214598 $T=167715 173875 0 0 $X=167315 $Y=173165
X89 2 VIA1_C_CDNS_724654214598 $T=167715 193895 0 0 $X=167315 $Y=193185
X90 13 VIA1_C_CDNS_724654214598 $T=168230 148400 0 0 $X=167830 $Y=147690
X91 2 VIA1_C_CDNS_724654214598 $T=168875 173875 0 0 $X=168475 $Y=173165
X92 2 VIA1_C_CDNS_724654214598 $T=168875 193895 0 0 $X=168475 $Y=193185
X93 4 VIA1_C_CDNS_724654214598 $T=169770 146620 0 0 $X=169370 $Y=145910
X94 14 VIA1_C_CDNS_724654214598 $T=170955 170315 0 0 $X=170555 $Y=169605
X95 15 VIA1_C_CDNS_724654214598 $T=170955 188555 0 0 $X=170555 $Y=187845
X96 13 VIA1_C_CDNS_724654214598 $T=171310 148400 0 0 $X=170910 $Y=147690
X97 2 VIA1_C_CDNS_724654214598 $T=172685 173875 0 0 $X=172285 $Y=173165
X98 2 VIA1_C_CDNS_724654214598 $T=172685 193895 0 0 $X=172285 $Y=193185
X99 4 VIA1_C_CDNS_724654214598 $T=172850 146620 0 0 $X=172450 $Y=145910
X100 15 VIA1_C_CDNS_724654214598 $T=174195 168535 0 0 $X=173795 $Y=167825
X101 13 VIA1_C_CDNS_724654214598 $T=174195 192115 0 0 $X=173795 $Y=191405
X102 13 VIA1_C_CDNS_724654214598 $T=174390 148400 0 0 $X=173990 $Y=147690
X103 2 VIA1_C_CDNS_724654214598 $T=175925 173875 0 0 $X=175525 $Y=173165
X104 2 VIA1_C_CDNS_724654214598 $T=175925 193895 0 0 $X=175525 $Y=193185
X105 4 VIA1_C_CDNS_724654214598 $T=175930 146620 0 0 $X=175530 $Y=145910
X106 13 VIA1_C_CDNS_724654214598 $T=177435 172095 0 0 $X=177035 $Y=171385
X107 14 VIA1_C_CDNS_724654214598 $T=177435 190335 0 0 $X=177035 $Y=189625
X108 13 VIA1_C_CDNS_724654214598 $T=177470 148400 0 0 $X=177070 $Y=147690
X109 4 VIA1_C_CDNS_724654214598 $T=179010 146620 0 0 $X=178610 $Y=145910
X110 2 VIA1_C_CDNS_724654214598 $T=179165 173875 0 0 $X=178765 $Y=173165
X111 2 VIA1_C_CDNS_724654214598 $T=179165 193895 0 0 $X=178765 $Y=193185
X112 13 VIA1_C_CDNS_724654214598 $T=180550 148400 0 0 $X=180150 $Y=147690
X113 14 VIA1_C_CDNS_724654214598 $T=180675 170315 0 0 $X=180275 $Y=169605
X114 15 VIA1_C_CDNS_724654214598 $T=180675 188555 0 0 $X=180275 $Y=187845
X115 2 VIA1_C_CDNS_724654214598 $T=182405 173875 0 0 $X=182005 $Y=173165
X116 2 VIA1_C_CDNS_724654214598 $T=182405 193895 0 0 $X=182005 $Y=193185
X117 13 VIA1_C_CDNS_724654214598 $T=183915 172095 0 0 $X=183515 $Y=171385
X118 15 VIA1_C_CDNS_724654214598 $T=183915 188555 0 0 $X=183515 $Y=187845
X119 2 VIA1_C_CDNS_724654214598 $T=185645 173875 0 0 $X=185245 $Y=173165
X120 2 VIA1_C_CDNS_724654214598 $T=185645 193895 0 0 $X=185245 $Y=193185
X121 15 VIA1_C_CDNS_724654214598 $T=187155 168535 0 0 $X=186755 $Y=167825
X122 13 VIA1_C_CDNS_724654214598 $T=187155 192115 0 0 $X=186755 $Y=191405
X123 2 VIA1_C_CDNS_724654214598 $T=188885 173875 0 0 $X=188485 $Y=173165
X124 2 VIA1_C_CDNS_724654214598 $T=188885 193895 0 0 $X=188485 $Y=193185
X125 14 VIA1_C_CDNS_724654214598 $T=189010 148400 0 0 $X=188610 $Y=147690
X126 13 VIA1_C_CDNS_724654214598 $T=190395 172095 0 0 $X=189995 $Y=171385
X127 14 VIA1_C_CDNS_724654214598 $T=190395 190335 0 0 $X=189995 $Y=189625
X128 6 VIA1_C_CDNS_724654214598 $T=190550 146620 0 0 $X=190150 $Y=145910
X129 14 VIA1_C_CDNS_724654214598 $T=192090 148400 0 0 $X=191690 $Y=147690
X130 2 VIA1_C_CDNS_724654214598 $T=192125 173875 0 0 $X=191725 $Y=173165
X131 2 VIA1_C_CDNS_724654214598 $T=192125 193895 0 0 $X=191725 $Y=193185
X132 6 VIA1_C_CDNS_724654214598 $T=193630 146620 0 0 $X=193230 $Y=145910
X133 14 VIA1_C_CDNS_724654214598 $T=193635 170315 0 0 $X=193235 $Y=169605
X134 13 VIA1_C_CDNS_724654214598 $T=193635 192115 0 0 $X=193235 $Y=191405
X135 14 VIA1_C_CDNS_724654214598 $T=195170 148400 0 0 $X=194770 $Y=147690
X136 2 VIA1_C_CDNS_724654214598 $T=195365 173875 0 0 $X=194965 $Y=173165
X137 2 VIA1_C_CDNS_724654214598 $T=195365 193895 0 0 $X=194965 $Y=193185
X138 6 VIA1_C_CDNS_724654214598 $T=196710 146620 0 0 $X=196310 $Y=145910
X139 13 VIA1_C_CDNS_724654214598 $T=196875 172095 0 0 $X=196475 $Y=171385
X140 15 VIA1_C_CDNS_724654214598 $T=196875 188555 0 0 $X=196475 $Y=187845
X141 14 VIA1_C_CDNS_724654214598 $T=198250 148400 0 0 $X=197850 $Y=147690
X142 2 VIA1_C_CDNS_724654214598 $T=198605 173875 0 0 $X=198205 $Y=173165
X143 2 VIA1_C_CDNS_724654214598 $T=198605 193895 0 0 $X=198205 $Y=193185
X144 6 VIA1_C_CDNS_724654214598 $T=199790 146620 0 0 $X=199390 $Y=145910
X145 15 VIA1_C_CDNS_724654214598 $T=200115 168535 0 0 $X=199715 $Y=167825
X146 13 VIA1_C_CDNS_724654214598 $T=200115 192115 0 0 $X=199715 $Y=191405
X147 14 VIA1_C_CDNS_724654214598 $T=201330 148400 0 0 $X=200930 $Y=147690
X148 2 VIA1_C_CDNS_724654214598 $T=201845 173875 0 0 $X=201445 $Y=173165
X149 2 VIA1_C_CDNS_724654214598 $T=201845 193895 0 0 $X=201445 $Y=193185
X150 6 VIA1_C_CDNS_724654214598 $T=202870 146620 0 0 $X=202470 $Y=145910
X151 13 VIA1_C_CDNS_724654214598 $T=203355 172095 0 0 $X=202955 $Y=171385
X152 14 VIA1_C_CDNS_724654214598 $T=203355 190335 0 0 $X=202955 $Y=189625
X153 14 VIA1_C_CDNS_724654214598 $T=204410 148400 0 0 $X=204010 $Y=147690
X154 2 VIA1_C_CDNS_724654214598 $T=205085 173875 0 0 $X=204685 $Y=173165
X155 2 VIA1_C_CDNS_724654214598 $T=205085 193895 0 0 $X=204685 $Y=193185
X156 14 VIA1_C_CDNS_724654214598 $T=206595 170315 0 0 $X=206195 $Y=169605
X157 13 VIA1_C_CDNS_724654214598 $T=206595 192115 0 0 $X=206195 $Y=191405
X158 2 VIA1_C_CDNS_724654214598 $T=208325 173875 0 0 $X=207925 $Y=173165
X159 2 VIA1_C_CDNS_724654214598 $T=208325 193895 0 0 $X=207925 $Y=193185
X160 14 VIA1_C_CDNS_724654214598 $T=209835 170315 0 0 $X=209435 $Y=169605
X161 15 VIA1_C_CDNS_724654214598 $T=209835 188555 0 0 $X=209435 $Y=187845
X162 2 VIA1_C_CDNS_724654214598 $T=211565 173875 0 0 $X=211165 $Y=173165
X163 2 VIA1_C_CDNS_724654214598 $T=211565 193895 0 0 $X=211165 $Y=193185
X164 15 VIA1_C_CDNS_724654214598 $T=212920 148400 0 0 $X=212520 $Y=147690
X165 15 VIA1_C_CDNS_724654214598 $T=213075 168535 0 0 $X=212675 $Y=167825
X166 13 VIA1_C_CDNS_724654214598 $T=213075 192115 0 0 $X=212675 $Y=191405
X167 5 VIA1_C_CDNS_724654214598 $T=214460 146620 0 0 $X=214060 $Y=145910
X168 2 VIA1_C_CDNS_724654214598 $T=214805 173875 0 0 $X=214405 $Y=173165
X169 2 VIA1_C_CDNS_724654214598 $T=214805 193895 0 0 $X=214405 $Y=193185
X170 15 VIA1_C_CDNS_724654214598 $T=216000 148400 0 0 $X=215600 $Y=147690
X171 13 VIA1_C_CDNS_724654214598 $T=216315 172095 0 0 $X=215915 $Y=171385
X172 14 VIA1_C_CDNS_724654214598 $T=216315 190335 0 0 $X=215915 $Y=189625
X173 5 VIA1_C_CDNS_724654214598 $T=217540 146620 0 0 $X=217140 $Y=145910
X174 2 VIA1_C_CDNS_724654214598 $T=218045 173875 0 0 $X=217645 $Y=173165
X175 2 VIA1_C_CDNS_724654214598 $T=218045 193895 0 0 $X=217645 $Y=193185
X176 15 VIA1_C_CDNS_724654214598 $T=219080 148400 0 0 $X=218680 $Y=147690
X177 14 VIA1_C_CDNS_724654214598 $T=219555 170315 0 0 $X=219155 $Y=169605
X178 15 VIA1_C_CDNS_724654214598 $T=219555 188555 0 0 $X=219155 $Y=187845
X179 5 VIA1_C_CDNS_724654214598 $T=220620 146620 0 0 $X=220220 $Y=145910
X180 2 VIA1_C_CDNS_724654214598 $T=221285 173875 0 0 $X=220885 $Y=173165
X181 2 VIA1_C_CDNS_724654214598 $T=221285 193895 0 0 $X=220885 $Y=193185
X182 2 VIA1_C_CDNS_724654214598 $T=221755 208575 0 0 $X=221355 $Y=207865
X183 15 VIA1_C_CDNS_724654214598 $T=222160 148400 0 0 $X=221760 $Y=147690
X184 2 VIA1_C_CDNS_724654214598 $T=223025 173875 0 0 $X=222625 $Y=173165
X185 2 VIA1_C_CDNS_724654214598 $T=223025 193895 0 0 $X=222625 $Y=193185
X186 5 VIA1_C_CDNS_724654214598 $T=223700 146620 0 0 $X=223300 $Y=145910
X187 15 VIA1_C_CDNS_724654214598 $T=225240 148400 0 0 $X=224840 $Y=147690
X188 5 VIA1_C_CDNS_724654214598 $T=226780 146620 0 0 $X=226380 $Y=145910
X189 15 VIA1_C_CDNS_724654214598 $T=228320 148400 0 0 $X=227920 $Y=147690
X190 8 VIA1_C_CDNS_724654214599 $T=162840 161880 0 0 $X=162440 $Y=161690
X191 8 VIA1_C_CDNS_724654214599 $T=164380 161880 0 0 $X=163980 $Y=161690
X192 8 VIA1_C_CDNS_724654214599 $T=165920 161880 0 0 $X=165520 $Y=161690
X193 8 VIA1_C_CDNS_724654214599 $T=167460 161880 0 0 $X=167060 $Y=161690
X194 8 VIA1_C_CDNS_724654214599 $T=169000 161880 0 0 $X=168600 $Y=161690
X195 8 VIA1_C_CDNS_724654214599 $T=170540 161880 0 0 $X=170140 $Y=161690
X196 8 VIA1_C_CDNS_724654214599 $T=172080 161880 0 0 $X=171680 $Y=161690
X197 8 VIA1_C_CDNS_724654214599 $T=173620 161880 0 0 $X=173220 $Y=161690
X198 8 VIA1_C_CDNS_724654214599 $T=175160 161880 0 0 $X=174760 $Y=161690
X199 8 VIA1_C_CDNS_724654214599 $T=176700 161880 0 0 $X=176300 $Y=161690
X200 8 VIA1_C_CDNS_724654214599 $T=178240 161880 0 0 $X=177840 $Y=161690
X201 8 VIA1_C_CDNS_724654214599 $T=179780 161880 0 0 $X=179380 $Y=161690
X202 8 VIA1_C_CDNS_724654214599 $T=189780 161880 0 0 $X=189380 $Y=161690
X203 8 VIA1_C_CDNS_724654214599 $T=191320 161880 0 0 $X=190920 $Y=161690
X204 8 VIA1_C_CDNS_724654214599 $T=192860 161880 0 0 $X=192460 $Y=161690
X205 8 VIA1_C_CDNS_724654214599 $T=194400 161880 0 0 $X=194000 $Y=161690
X206 8 VIA1_C_CDNS_724654214599 $T=195940 161880 0 0 $X=195540 $Y=161690
X207 8 VIA1_C_CDNS_724654214599 $T=197480 161880 0 0 $X=197080 $Y=161690
X208 8 VIA1_C_CDNS_724654214599 $T=199020 161880 0 0 $X=198620 $Y=161690
X209 8 VIA1_C_CDNS_724654214599 $T=200560 161880 0 0 $X=200160 $Y=161690
X210 8 VIA1_C_CDNS_724654214599 $T=202100 161880 0 0 $X=201700 $Y=161690
X211 8 VIA1_C_CDNS_724654214599 $T=203640 161880 0 0 $X=203240 $Y=161690
X212 8 VIA1_C_CDNS_724654214599 $T=213690 161880 0 0 $X=213290 $Y=161690
X213 8 VIA1_C_CDNS_724654214599 $T=215230 161880 0 0 $X=214830 $Y=161690
X214 8 VIA1_C_CDNS_724654214599 $T=216770 161880 0 0 $X=216370 $Y=161690
X215 8 VIA1_C_CDNS_724654214599 $T=218310 161880 0 0 $X=217910 $Y=161690
X216 8 VIA1_C_CDNS_724654214599 $T=219850 161880 0 0 $X=219450 $Y=161690
X217 8 VIA1_C_CDNS_724654214599 $T=221390 161880 0 0 $X=220990 $Y=161690
X218 8 VIA1_C_CDNS_724654214599 $T=222930 161880 0 0 $X=222530 $Y=161690
X219 8 VIA1_C_CDNS_724654214599 $T=224470 161880 0 0 $X=224070 $Y=161690
X220 8 VIA1_C_CDNS_724654214599 $T=226010 161880 0 0 $X=225610 $Y=161690
X221 8 VIA1_C_CDNS_724654214599 $T=227550 161880 0 0 $X=227150 $Y=161690
X222 3 VIA1_C_CDNS_7246542145910 $T=18545 65405 0 0 $X=18355 $Y=65215
X223 3 VIA1_C_CDNS_7246542145910 $T=21085 65405 0 0 $X=20895 $Y=65215
X224 3 VIA1_C_CDNS_7246542145910 $T=23625 65405 0 0 $X=23435 $Y=65215
X225 3 VIA1_C_CDNS_7246542145910 $T=26165 65405 0 0 $X=25975 $Y=65215
X226 3 VIA1_C_CDNS_7246542145910 $T=28705 65405 0 0 $X=28515 $Y=65215
X227 3 VIA1_C_CDNS_7246542145910 $T=31245 65405 0 0 $X=31055 $Y=65215
X228 3 VIA1_C_CDNS_7246542145910 $T=33785 65405 0 0 $X=33595 $Y=65215
X229 3 VIA1_C_CDNS_7246542145910 $T=36325 65405 0 0 $X=36135 $Y=65215
X230 3 VIA1_C_CDNS_7246542145911 $T=43480 65295 0 0 $X=42560 $Y=65105
X231 3 VIA1_C_CDNS_7246542145911 $T=46020 65295 0 0 $X=45100 $Y=65105
X232 3 VIA1_C_CDNS_7246542145911 $T=48560 65295 0 0 $X=47640 $Y=65105
X233 3 VIA1_C_CDNS_7246542145911 $T=51100 65295 0 0 $X=50180 $Y=65105
X234 3 VIA1_C_CDNS_7246542145911 $T=53640 65295 0 0 $X=52720 $Y=65105
X235 3 VIA1_C_CDNS_7246542145911 $T=56180 65295 0 0 $X=55260 $Y=65105
X236 3 VIA1_C_CDNS_7246542145911 $T=58720 65295 0 0 $X=57800 $Y=65105
X237 3 VIA1_C_CDNS_7246542145911 $T=61260 65295 0 0 $X=60340 $Y=65105
X238 12 VIA1_C_CDNS_7246542145911 $T=139060 201685 0 0 $X=138140 $Y=201495
X239 12 VIA1_C_CDNS_7246542145911 $T=141600 201685 0 0 $X=140680 $Y=201495
X240 8 VIA1_C_CDNS_7246542145911 $T=148620 201685 0 0 $X=147700 $Y=201495
X241 8 VIA1_C_CDNS_7246542145911 $T=151160 201685 0 0 $X=150240 $Y=201495
X242 2 VIA1_C_CDNS_7246542145912 $T=22280 170260 0 0 $X=22140 $Y=169550
X243 2 VIA1_C_CDNS_7246542145912 $T=22980 170260 0 0 $X=22840 $Y=169550
X244 2 VIA1_C_CDNS_7246542145912 $T=22980 187940 0 0 $X=22840 $Y=187230
X245 16 VIA1_C_CDNS_7246542145912 $T=33520 166700 0 0 $X=33380 $Y=165990
X246 17 VIA1_C_CDNS_7246542145912 $T=33520 186160 0 0 $X=33380 $Y=185450
X247 2 VIA1_C_CDNS_7246542145912 $T=34220 170260 0 0 $X=34080 $Y=169550
X248 2 VIA1_C_CDNS_7246542145912 $T=34220 187940 0 0 $X=34080 $Y=187230
X249 17 VIA1_C_CDNS_7246542145912 $T=44760 168480 0 0 $X=44620 $Y=167770
X250 16 VIA1_C_CDNS_7246542145912 $T=44760 184380 0 0 $X=44620 $Y=183670
X251 2 VIA1_C_CDNS_7246542145912 $T=45460 170260 0 0 $X=45320 $Y=169550
X252 2 VIA1_C_CDNS_7246542145912 $T=45460 187940 0 0 $X=45320 $Y=187230
X253 16 VIA1_C_CDNS_7246542145912 $T=56000 166700 0 0 $X=55860 $Y=165990
X254 17 VIA1_C_CDNS_7246542145912 $T=56000 186160 0 0 $X=55860 $Y=185450
X255 2 VIA1_C_CDNS_7246542145912 $T=56700 170260 0 0 $X=56560 $Y=169550
X256 2 VIA1_C_CDNS_7246542145912 $T=56700 187940 0 0 $X=56560 $Y=187230
X257 17 VIA1_C_CDNS_7246542145912 $T=67240 168480 0 0 $X=67100 $Y=167770
X258 16 VIA1_C_CDNS_7246542145912 $T=67240 184380 0 0 $X=67100 $Y=183670
X259 2 VIA1_C_CDNS_7246542145912 $T=67940 170260 0 0 $X=67800 $Y=169550
X260 2 VIA1_C_CDNS_7246542145912 $T=67940 187940 0 0 $X=67800 $Y=187230
X261 16 VIA1_C_CDNS_7246542145912 $T=78480 166700 0 0 $X=78340 $Y=165990
X262 17 VIA1_C_CDNS_7246542145912 $T=78480 186160 0 0 $X=78340 $Y=185450
X263 2 VIA1_C_CDNS_7246542145912 $T=79180 170260 0 0 $X=79040 $Y=169550
X264 2 VIA1_C_CDNS_7246542145912 $T=79180 187940 0 0 $X=79040 $Y=187230
X265 17 VIA1_C_CDNS_7246542145912 $T=89720 168480 0 0 $X=89580 $Y=167770
X266 16 VIA1_C_CDNS_7246542145912 $T=89720 184380 0 0 $X=89580 $Y=183670
X267 2 VIA1_C_CDNS_7246542145912 $T=90420 170260 0 0 $X=90280 $Y=169550
X268 2 VIA1_C_CDNS_7246542145912 $T=90420 187940 0 0 $X=90280 $Y=187230
X269 16 VIA1_C_CDNS_7246542145912 $T=100960 166700 0 0 $X=100820 $Y=165990
X270 17 VIA1_C_CDNS_7246542145912 $T=100960 186160 0 0 $X=100820 $Y=185450
X271 2 VIA1_C_CDNS_7246542145912 $T=101660 170260 0 0 $X=101520 $Y=169550
X272 2 VIA1_C_CDNS_7246542145912 $T=101660 187940 0 0 $X=101520 $Y=187230
X273 17 VIA1_C_CDNS_7246542145912 $T=112200 168480 0 0 $X=112060 $Y=167770
X274 16 VIA1_C_CDNS_7246542145912 $T=112200 184380 0 0 $X=112060 $Y=183670
X275 2 VIA1_C_CDNS_7246542145912 $T=112900 170260 0 0 $X=112760 $Y=169550
X276 2 VIA1_C_CDNS_7246542145912 $T=112900 187940 0 0 $X=112760 $Y=187230
X277 16 VIA2_C_CDNS_7246542145913 $T=7190 201560 0 0 $X=6480 $Y=201420
X278 16 VIA1_C_CDNS_7246542145914 $T=28250 201560 0 0 $X=27590 $Y=201370
X279 16 VIA1_C_CDNS_7246542145914 $T=39490 201560 0 0 $X=38830 $Y=201370
X280 16 VIA1_C_CDNS_7246542145914 $T=50730 201560 0 0 $X=50070 $Y=201370
X281 16 VIA1_C_CDNS_7246542145914 $T=61970 201560 0 0 $X=61310 $Y=201370
X282 16 VIA1_C_CDNS_7246542145914 $T=73210 201560 0 0 $X=72550 $Y=201370
X283 16 VIA1_C_CDNS_7246542145914 $T=84450 201560 0 0 $X=83790 $Y=201370
X284 16 VIA1_C_CDNS_7246542145914 $T=95690 201560 0 0 $X=95030 $Y=201370
X285 16 VIA1_C_CDNS_7246542145914 $T=106930 201560 0 0 $X=106270 $Y=201370
X286 17 VIA1_C_CDNS_7246542145915 $T=169915 187385 0 0 $X=168945 $Y=187195
X287 17 VIA1_C_CDNS_7246542145915 $T=169915 207405 0 0 $X=168945 $Y=207215
X288 17 VIA1_C_CDNS_7246542145915 $T=173155 187385 0 0 $X=172185 $Y=187195
X289 17 VIA1_C_CDNS_7246542145915 $T=173155 207405 0 0 $X=172185 $Y=207215
X290 17 VIA1_C_CDNS_7246542145915 $T=176395 187385 0 0 $X=175425 $Y=187195
X291 17 VIA1_C_CDNS_7246542145915 $T=176395 207405 0 0 $X=175425 $Y=207215
X292 17 VIA1_C_CDNS_7246542145915 $T=179635 187385 0 0 $X=178665 $Y=187195
X293 17 VIA1_C_CDNS_7246542145915 $T=179635 207405 0 0 $X=178665 $Y=207215
X294 17 VIA1_C_CDNS_7246542145915 $T=182875 187385 0 0 $X=181905 $Y=187195
X295 17 VIA1_C_CDNS_7246542145915 $T=182875 207405 0 0 $X=181905 $Y=207215
X296 17 VIA1_C_CDNS_7246542145915 $T=186115 187385 0 0 $X=185145 $Y=187195
X297 17 VIA1_C_CDNS_7246542145915 $T=186115 207405 0 0 $X=185145 $Y=207215
X298 17 VIA1_C_CDNS_7246542145915 $T=189355 187385 0 0 $X=188385 $Y=187195
X299 17 VIA1_C_CDNS_7246542145915 $T=189355 207405 0 0 $X=188385 $Y=207215
X300 17 VIA1_C_CDNS_7246542145915 $T=192595 187385 0 0 $X=191625 $Y=187195
X301 17 VIA1_C_CDNS_7246542145915 $T=192595 207405 0 0 $X=191625 $Y=207215
X302 17 VIA1_C_CDNS_7246542145915 $T=195835 187385 0 0 $X=194865 $Y=187195
X303 17 VIA1_C_CDNS_7246542145915 $T=195835 207405 0 0 $X=194865 $Y=207215
X304 17 VIA1_C_CDNS_7246542145915 $T=199075 187385 0 0 $X=198105 $Y=187195
X305 17 VIA1_C_CDNS_7246542145915 $T=199075 207405 0 0 $X=198105 $Y=207215
X306 17 VIA1_C_CDNS_7246542145915 $T=202315 187385 0 0 $X=201345 $Y=187195
X307 17 VIA1_C_CDNS_7246542145915 $T=202315 207405 0 0 $X=201345 $Y=207215
X308 17 VIA1_C_CDNS_7246542145915 $T=205555 187385 0 0 $X=204585 $Y=187195
X309 17 VIA1_C_CDNS_7246542145915 $T=205555 207405 0 0 $X=204585 $Y=207215
X310 17 VIA1_C_CDNS_7246542145915 $T=208795 187385 0 0 $X=207825 $Y=187195
X311 17 VIA1_C_CDNS_7246542145915 $T=208795 207405 0 0 $X=207825 $Y=207215
X312 17 VIA1_C_CDNS_7246542145915 $T=212035 187385 0 0 $X=211065 $Y=187195
X313 17 VIA1_C_CDNS_7246542145915 $T=212035 207405 0 0 $X=211065 $Y=207215
X314 17 VIA1_C_CDNS_7246542145915 $T=215275 187385 0 0 $X=214305 $Y=187195
X315 17 VIA1_C_CDNS_7246542145915 $T=215275 207405 0 0 $X=214305 $Y=207215
X316 17 VIA1_C_CDNS_7246542145915 $T=218515 187385 0 0 $X=217545 $Y=187195
X317 17 VIA1_C_CDNS_7246542145915 $T=218515 207405 0 0 $X=217545 $Y=207215
X318 2 VIA1_C_CDNS_7246542145916 $T=11740 170260 0 0 $X=11550 $Y=169600
X319 2 VIA1_C_CDNS_7246542145916 $T=11740 187940 0 0 $X=11550 $Y=187280
X320 2 VIA1_C_CDNS_7246542145916 $T=17010 187940 0 0 $X=16820 $Y=187280
X321 2 VIA1_C_CDNS_7246542145916 $T=22280 187940 0 0 $X=22090 $Y=187280
X322 16 VIA1_C_CDNS_7246542145916 $T=28250 184380 0 0 $X=28060 $Y=183720
X323 16 VIA1_C_CDNS_7246542145916 $T=39490 184380 0 0 $X=39300 $Y=183720
X324 16 VIA1_C_CDNS_7246542145916 $T=50730 184380 0 0 $X=50540 $Y=183720
X325 16 VIA1_C_CDNS_7246542145916 $T=61970 184380 0 0 $X=61780 $Y=183720
X326 16 VIA1_C_CDNS_7246542145916 $T=73210 184380 0 0 $X=73020 $Y=183720
X327 16 VIA1_C_CDNS_7246542145916 $T=84450 184380 0 0 $X=84260 $Y=183720
X328 16 VIA1_C_CDNS_7246542145916 $T=95690 184380 0 0 $X=95500 $Y=183720
X329 16 VIA1_C_CDNS_7246542145916 $T=106930 184380 0 0 $X=106740 $Y=183720
X330 2 VIA1_C_CDNS_7246542145916 $T=118170 187940 0 0 $X=117980 $Y=187280
X331 2 VIA1_C_CDNS_7246542145916 $T=123440 170260 0 0 $X=123250 $Y=169600
X332 2 VIA1_C_CDNS_7246542145916 $T=123440 187940 0 0 $X=123250 $Y=187280
X333 1 VIA2_C_CDNS_7246542145917 $T=15905 4500 0 0 $X=13335 $Y=3230
X334 1 VIA2_C_CDNS_7246542145917 $T=62500 4500 0 0 $X=59930 $Y=3230
X335 2 VIA2_C_CDNS_7246542145918 $T=9220 170260 0 0 $X=8250 $Y=169600
X336 2 VIA2_C_CDNS_7246542145918 $T=9220 187940 0 0 $X=8250 $Y=187280
X337 2 VIA2_C_CDNS_7246542145918 $T=125960 170260 0 0 $X=124990 $Y=169600
X338 2 VIA2_C_CDNS_7246542145918 $T=125960 187940 0 0 $X=124990 $Y=187280
X339 2 VIA2_C_CDNS_7246542145918 $T=162885 173875 0 0 $X=161915 $Y=173215
X340 2 VIA2_C_CDNS_7246542145918 $T=162885 193895 0 0 $X=161915 $Y=193235
X341 2 VIA2_C_CDNS_7246542145918 $T=162885 208575 0 0 $X=161915 $Y=207915
X342 2 VIA2_C_CDNS_7246542145918 $T=225545 173875 0 0 $X=224575 $Y=173215
X343 2 VIA2_C_CDNS_7246542145918 $T=225545 193895 0 0 $X=224575 $Y=193235
X344 2 VIA2_C_CDNS_7246542145918 $T=225545 208575 0 0 $X=224575 $Y=207915
X345 16 VIA2_C_CDNS_7246542145919 $T=7190 166700 0 0 $X=6480 $Y=166040
X346 16 VIA2_C_CDNS_7246542145919 $T=7190 184380 0 0 $X=6480 $Y=183720
X347 17 VIA2_C_CDNS_7246542145919 $T=127990 168480 0 0 $X=127280 $Y=167820
X348 17 VIA2_C_CDNS_7246542145919 $T=127990 186160 0 0 $X=127280 $Y=185500
X349 13 VIA2_C_CDNS_7246542145919 $T=160855 172095 0 0 $X=160145 $Y=171435
X350 13 VIA2_C_CDNS_7246542145919 $T=160855 192115 0 0 $X=160145 $Y=191455
X351 14 VIA2_C_CDNS_7246542145919 $T=227575 170315 0 0 $X=226865 $Y=169655
X352 14 VIA2_C_CDNS_7246542145919 $T=227575 190335 0 0 $X=226865 $Y=189675
X353 15 VIA2_C_CDNS_7246542145919 $T=229355 168535 0 0 $X=228645 $Y=167875
X354 15 VIA2_C_CDNS_7246542145919 $T=229355 188555 0 0 $X=228645 $Y=187895
X355 1 VIA1_C_CDNS_7246542145920 $T=117240 7840 0 90 $X=116270 $Y=7440
X356 1 VIA1_C_CDNS_7246542145920 $T=117240 38150 0 90 $X=116270 $Y=37750
X357 1 VIA1_C_CDNS_7246542145920 $T=117240 39310 0 90 $X=116270 $Y=38910
X358 1 VIA1_C_CDNS_7246542145920 $T=117240 69390 0 90 $X=116270 $Y=68990
X359 1 VIA1_C_CDNS_7246542145920 $T=117240 70550 0 90 $X=116270 $Y=70150
X360 1 VIA1_C_CDNS_7246542145920 $T=117240 100860 0 90 $X=116270 $Y=100460
X361 1 VIA1_C_CDNS_7246542145920 $T=154205 7780 0 90 $X=153235 $Y=7380
X362 1 VIA1_C_CDNS_7246542145920 $T=154205 38090 0 90 $X=153235 $Y=37690
X363 1 VIA1_C_CDNS_7246542145920 $T=154205 39250 0 90 $X=153235 $Y=38850
X364 1 VIA1_C_CDNS_7246542145920 $T=154205 69330 0 90 $X=153235 $Y=68930
X365 1 VIA1_C_CDNS_7246542145920 $T=154205 70490 0 90 $X=153235 $Y=70090
X366 1 VIA1_C_CDNS_7246542145920 $T=154205 100800 0 90 $X=153235 $Y=100400
X367 5 VIA1_C_CDNS_7246542145921 $T=83930 23110 0 90 $X=83220 $Y=22450
X368 5 VIA1_C_CDNS_7246542145921 $T=83930 54350 0 90 $X=83220 $Y=53690
X369 5 VIA1_C_CDNS_7246542145921 $T=83930 85590 0 90 $X=83220 $Y=84930
X370 6 VIA1_C_CDNS_7246542145921 $T=120895 23050 0 90 $X=120185 $Y=22390
X371 6 VIA1_C_CDNS_7246542145921 $T=120895 54290 0 90 $X=120185 $Y=53630
X372 6 VIA1_C_CDNS_7246542145921 $T=120895 85530 0 90 $X=120185 $Y=84870
X373 4 VIA2_C_CDNS_7246542145922 $T=17790 130490 0 0 $X=17650 $Y=130300
X374 7 VIA2_C_CDNS_7246542145922 $T=17790 131270 0 0 $X=17650 $Y=131080
X375 4 VIA2_C_CDNS_7246542145922 $T=20880 130490 0 0 $X=20740 $Y=130300
X376 7 VIA2_C_CDNS_7246542145922 $T=21500 131270 0 0 $X=21360 $Y=131080
X377 4 VIA2_C_CDNS_7246542145922 $T=24590 130490 0 0 $X=24450 $Y=130300
X378 7 VIA2_C_CDNS_7246542145922 $T=24590 131270 0 0 $X=24450 $Y=131080
X379 4 VIA2_C_CDNS_7246542145922 $T=27680 130490 0 0 $X=27540 $Y=130300
X380 7 VIA2_C_CDNS_7246542145922 $T=28300 131270 0 0 $X=28160 $Y=131080
X381 4 VIA2_C_CDNS_7246542145922 $T=31390 130490 0 0 $X=31250 $Y=130300
X382 7 VIA2_C_CDNS_7246542145922 $T=31390 131270 0 0 $X=31250 $Y=131080
X383 4 VIA2_C_CDNS_7246542145922 $T=34480 130490 0 0 $X=34340 $Y=130300
X384 7 VIA2_C_CDNS_7246542145922 $T=35100 131270 0 0 $X=34960 $Y=131080
X385 4 VIA2_C_CDNS_7246542145922 $T=38190 130490 0 0 $X=38050 $Y=130300
X386 7 VIA2_C_CDNS_7246542145922 $T=38190 131270 0 0 $X=38050 $Y=131080
X387 4 VIA2_C_CDNS_7246542145922 $T=41280 130490 0 0 $X=41140 $Y=130300
X388 7 VIA2_C_CDNS_7246542145922 $T=41900 131270 0 0 $X=41760 $Y=131080
X389 4 VIA2_C_CDNS_7246542145922 $T=44990 130490 0 0 $X=44850 $Y=130300
X390 7 VIA2_C_CDNS_7246542145922 $T=44990 131270 0 0 $X=44850 $Y=131080
X391 4 VIA2_C_CDNS_7246542145922 $T=48080 130490 0 0 $X=47940 $Y=130300
X392 7 VIA2_C_CDNS_7246542145922 $T=48700 131270 0 0 $X=48560 $Y=131080
X393 4 VIA2_C_CDNS_7246542145922 $T=51790 130490 0 0 $X=51650 $Y=130300
X394 7 VIA2_C_CDNS_7246542145922 $T=51790 131270 0 0 $X=51650 $Y=131080
X395 4 VIA2_C_CDNS_7246542145922 $T=54880 130490 0 0 $X=54740 $Y=130300
X396 7 VIA2_C_CDNS_7246542145922 $T=55500 131270 0 0 $X=55360 $Y=131080
X397 4 VIA2_C_CDNS_7246542145922 $T=58590 130490 0 0 $X=58450 $Y=130300
X398 7 VIA2_C_CDNS_7246542145922 $T=58590 131270 0 0 $X=58450 $Y=131080
X399 4 VIA2_C_CDNS_7246542145922 $T=61680 130490 0 0 $X=61540 $Y=130300
X400 7 VIA2_C_CDNS_7246542145922 $T=62300 131270 0 0 $X=62160 $Y=131080
X401 11 VIA1_C_CDNS_7246542145923 $T=14390 117740 0 0 $X=13680 $Y=117600
X402 11 VIA1_C_CDNS_7246542145923 $T=14390 144020 0 0 $X=13680 $Y=143880
X403 11 VIA1_C_CDNS_7246542145923 $T=17790 117740 0 0 $X=17080 $Y=117600
X404 11 VIA1_C_CDNS_7246542145923 $T=17790 144020 0 0 $X=17080 $Y=143880
X405 11 VIA1_C_CDNS_7246542145923 $T=21190 117740 0 0 $X=20480 $Y=117600
X406 11 VIA1_C_CDNS_7246542145923 $T=21190 144020 0 0 $X=20480 $Y=143880
X407 11 VIA1_C_CDNS_7246542145923 $T=24590 117740 0 0 $X=23880 $Y=117600
X408 11 VIA1_C_CDNS_7246542145923 $T=24590 144020 0 0 $X=23880 $Y=143880
X409 11 VIA1_C_CDNS_7246542145923 $T=27990 117740 0 0 $X=27280 $Y=117600
X410 11 VIA1_C_CDNS_7246542145923 $T=27990 144020 0 0 $X=27280 $Y=143880
X411 11 VIA1_C_CDNS_7246542145923 $T=31390 117740 0 0 $X=30680 $Y=117600
X412 11 VIA1_C_CDNS_7246542145923 $T=31390 144020 0 0 $X=30680 $Y=143880
X413 11 VIA1_C_CDNS_7246542145923 $T=34790 117740 0 0 $X=34080 $Y=117600
X414 11 VIA1_C_CDNS_7246542145923 $T=34790 144020 0 0 $X=34080 $Y=143880
X415 11 VIA1_C_CDNS_7246542145923 $T=38190 117740 0 0 $X=37480 $Y=117600
X416 11 VIA1_C_CDNS_7246542145923 $T=38190 144020 0 0 $X=37480 $Y=143880
X417 11 VIA1_C_CDNS_7246542145923 $T=41590 117740 0 0 $X=40880 $Y=117600
X418 11 VIA1_C_CDNS_7246542145923 $T=41590 144020 0 0 $X=40880 $Y=143880
X419 11 VIA1_C_CDNS_7246542145923 $T=44990 117740 0 0 $X=44280 $Y=117600
X420 11 VIA1_C_CDNS_7246542145923 $T=44990 144020 0 0 $X=44280 $Y=143880
X421 11 VIA1_C_CDNS_7246542145923 $T=48390 117740 0 0 $X=47680 $Y=117600
X422 11 VIA1_C_CDNS_7246542145923 $T=48390 144020 0 0 $X=47680 $Y=143880
X423 11 VIA1_C_CDNS_7246542145923 $T=51790 117740 0 0 $X=51080 $Y=117600
X424 11 VIA1_C_CDNS_7246542145923 $T=51790 144020 0 0 $X=51080 $Y=143880
X425 11 VIA1_C_CDNS_7246542145923 $T=55190 117740 0 0 $X=54480 $Y=117600
X426 11 VIA1_C_CDNS_7246542145923 $T=55190 144020 0 0 $X=54480 $Y=143880
X427 11 VIA1_C_CDNS_7246542145923 $T=58590 117740 0 0 $X=57880 $Y=117600
X428 11 VIA1_C_CDNS_7246542145923 $T=58590 144020 0 0 $X=57880 $Y=143880
X429 11 VIA1_C_CDNS_7246542145923 $T=61990 117740 0 0 $X=61280 $Y=117600
X430 11 VIA1_C_CDNS_7246542145923 $T=61990 144020 0 0 $X=61280 $Y=143880
X431 11 VIA1_C_CDNS_7246542145923 $T=65390 117740 0 0 $X=64680 $Y=117600
X432 11 VIA1_C_CDNS_7246542145923 $T=65390 144020 0 0 $X=64680 $Y=143880
X433 11 VIA2_C_CDNS_7246542145924 $T=13120 115960 0 0 $X=12980 $Y=115250
X434 11 VIA2_C_CDNS_7246542145924 $T=13120 145800 0 0 $X=12980 $Y=145090
X435 11 VIA2_C_CDNS_7246542145924 $T=14390 115960 0 0 $X=14250 $Y=115250
X436 11 VIA2_C_CDNS_7246542145924 $T=14390 145800 0 0 $X=14250 $Y=145090
X437 11 VIA2_C_CDNS_7246542145924 $T=15660 115960 0 0 $X=15520 $Y=115250
X438 11 VIA2_C_CDNS_7246542145924 $T=15660 145800 0 0 $X=15520 $Y=145090
X439 11 VIA2_C_CDNS_7246542145924 $T=16520 115960 0 0 $X=16380 $Y=115250
X440 11 VIA2_C_CDNS_7246542145924 $T=16520 145800 0 0 $X=16380 $Y=145090
X441 11 VIA2_C_CDNS_7246542145924 $T=17790 115960 0 0 $X=17650 $Y=115250
X442 11 VIA2_C_CDNS_7246542145924 $T=17790 145800 0 0 $X=17650 $Y=145090
X443 16 VIA2_C_CDNS_7246542145924 $T=19060 112400 0 0 $X=18920 $Y=111690
X444 17 VIA2_C_CDNS_7246542145924 $T=19060 149360 0 0 $X=18920 $Y=148650
X445 11 VIA2_C_CDNS_7246542145924 $T=19920 115960 0 0 $X=19780 $Y=115250
X446 11 VIA2_C_CDNS_7246542145924 $T=19920 145800 0 0 $X=19780 $Y=145090
X447 11 VIA2_C_CDNS_7246542145924 $T=21190 115960 0 0 $X=21050 $Y=115250
X448 11 VIA2_C_CDNS_7246542145924 $T=21190 145800 0 0 $X=21050 $Y=145090
X449 17 VIA2_C_CDNS_7246542145924 $T=22460 114180 0 0 $X=22320 $Y=113470
X450 16 VIA2_C_CDNS_7246542145924 $T=22460 147580 0 0 $X=22320 $Y=146870
X451 11 VIA2_C_CDNS_7246542145924 $T=23320 115960 0 0 $X=23180 $Y=115250
X452 11 VIA2_C_CDNS_7246542145924 $T=23320 145800 0 0 $X=23180 $Y=145090
X453 11 VIA2_C_CDNS_7246542145924 $T=24590 115960 0 0 $X=24450 $Y=115250
X454 11 VIA2_C_CDNS_7246542145924 $T=24590 145800 0 0 $X=24450 $Y=145090
X455 16 VIA2_C_CDNS_7246542145924 $T=25860 112400 0 0 $X=25720 $Y=111690
X456 17 VIA2_C_CDNS_7246542145924 $T=25860 149360 0 0 $X=25720 $Y=148650
X457 11 VIA2_C_CDNS_7246542145924 $T=26720 115960 0 0 $X=26580 $Y=115250
X458 11 VIA2_C_CDNS_7246542145924 $T=26720 145800 0 0 $X=26580 $Y=145090
X459 11 VIA2_C_CDNS_7246542145924 $T=27990 115960 0 0 $X=27850 $Y=115250
X460 11 VIA2_C_CDNS_7246542145924 $T=27990 145800 0 0 $X=27850 $Y=145090
X461 17 VIA2_C_CDNS_7246542145924 $T=29260 114180 0 0 $X=29120 $Y=113470
X462 16 VIA2_C_CDNS_7246542145924 $T=29260 147580 0 0 $X=29120 $Y=146870
X463 11 VIA2_C_CDNS_7246542145924 $T=30120 115960 0 0 $X=29980 $Y=115250
X464 11 VIA2_C_CDNS_7246542145924 $T=30120 145800 0 0 $X=29980 $Y=145090
X465 11 VIA2_C_CDNS_7246542145924 $T=31390 115960 0 0 $X=31250 $Y=115250
X466 11 VIA2_C_CDNS_7246542145924 $T=31390 145800 0 0 $X=31250 $Y=145090
X467 16 VIA2_C_CDNS_7246542145924 $T=32660 112400 0 0 $X=32520 $Y=111690
X468 17 VIA2_C_CDNS_7246542145924 $T=32660 149360 0 0 $X=32520 $Y=148650
X469 11 VIA2_C_CDNS_7246542145924 $T=33520 115960 0 0 $X=33380 $Y=115250
X470 11 VIA2_C_CDNS_7246542145924 $T=33520 145800 0 0 $X=33380 $Y=145090
X471 11 VIA2_C_CDNS_7246542145924 $T=34790 115960 0 0 $X=34650 $Y=115250
X472 11 VIA2_C_CDNS_7246542145924 $T=34790 145800 0 0 $X=34650 $Y=145090
X473 17 VIA2_C_CDNS_7246542145924 $T=36060 114180 0 0 $X=35920 $Y=113470
X474 16 VIA2_C_CDNS_7246542145924 $T=36060 147580 0 0 $X=35920 $Y=146870
X475 11 VIA2_C_CDNS_7246542145924 $T=36920 115960 0 0 $X=36780 $Y=115250
X476 11 VIA2_C_CDNS_7246542145924 $T=36920 145800 0 0 $X=36780 $Y=145090
X477 11 VIA2_C_CDNS_7246542145924 $T=38190 115960 0 0 $X=38050 $Y=115250
X478 11 VIA2_C_CDNS_7246542145924 $T=38190 145800 0 0 $X=38050 $Y=145090
X479 16 VIA2_C_CDNS_7246542145924 $T=39460 112400 0 0 $X=39320 $Y=111690
X480 17 VIA2_C_CDNS_7246542145924 $T=39460 149360 0 0 $X=39320 $Y=148650
X481 11 VIA2_C_CDNS_7246542145924 $T=40320 115960 0 0 $X=40180 $Y=115250
X482 11 VIA2_C_CDNS_7246542145924 $T=40320 145800 0 0 $X=40180 $Y=145090
X483 11 VIA2_C_CDNS_7246542145924 $T=41590 115960 0 0 $X=41450 $Y=115250
X484 11 VIA2_C_CDNS_7246542145924 $T=41590 145800 0 0 $X=41450 $Y=145090
X485 17 VIA2_C_CDNS_7246542145924 $T=42860 114180 0 0 $X=42720 $Y=113470
X486 16 VIA2_C_CDNS_7246542145924 $T=42860 147580 0 0 $X=42720 $Y=146870
X487 11 VIA2_C_CDNS_7246542145924 $T=43720 115960 0 0 $X=43580 $Y=115250
X488 11 VIA2_C_CDNS_7246542145924 $T=43720 145800 0 0 $X=43580 $Y=145090
X489 11 VIA2_C_CDNS_7246542145924 $T=44990 115960 0 0 $X=44850 $Y=115250
X490 11 VIA2_C_CDNS_7246542145924 $T=44990 145800 0 0 $X=44850 $Y=145090
X491 16 VIA2_C_CDNS_7246542145924 $T=46260 112400 0 0 $X=46120 $Y=111690
X492 17 VIA2_C_CDNS_7246542145924 $T=46260 149360 0 0 $X=46120 $Y=148650
X493 11 VIA2_C_CDNS_7246542145924 $T=47120 115960 0 0 $X=46980 $Y=115250
X494 11 VIA2_C_CDNS_7246542145924 $T=47120 145800 0 0 $X=46980 $Y=145090
X495 11 VIA2_C_CDNS_7246542145924 $T=48390 115960 0 0 $X=48250 $Y=115250
X496 11 VIA2_C_CDNS_7246542145924 $T=48390 145800 0 0 $X=48250 $Y=145090
X497 17 VIA2_C_CDNS_7246542145924 $T=49660 114180 0 0 $X=49520 $Y=113470
X498 16 VIA2_C_CDNS_7246542145924 $T=49660 147580 0 0 $X=49520 $Y=146870
X499 11 VIA2_C_CDNS_7246542145924 $T=50520 115960 0 0 $X=50380 $Y=115250
X500 11 VIA2_C_CDNS_7246542145924 $T=50520 145800 0 0 $X=50380 $Y=145090
X501 11 VIA2_C_CDNS_7246542145924 $T=51790 115960 0 0 $X=51650 $Y=115250
X502 11 VIA2_C_CDNS_7246542145924 $T=51790 145800 0 0 $X=51650 $Y=145090
X503 16 VIA2_C_CDNS_7246542145924 $T=53060 112400 0 0 $X=52920 $Y=111690
X504 17 VIA2_C_CDNS_7246542145924 $T=53060 149360 0 0 $X=52920 $Y=148650
X505 11 VIA2_C_CDNS_7246542145924 $T=53920 115960 0 0 $X=53780 $Y=115250
X506 11 VIA2_C_CDNS_7246542145924 $T=53920 145800 0 0 $X=53780 $Y=145090
X507 11 VIA2_C_CDNS_7246542145924 $T=55190 115960 0 0 $X=55050 $Y=115250
X508 11 VIA2_C_CDNS_7246542145924 $T=55190 145800 0 0 $X=55050 $Y=145090
X509 17 VIA2_C_CDNS_7246542145924 $T=56460 114180 0 0 $X=56320 $Y=113470
X510 16 VIA2_C_CDNS_7246542145924 $T=56460 147580 0 0 $X=56320 $Y=146870
X511 11 VIA2_C_CDNS_7246542145924 $T=57320 115960 0 0 $X=57180 $Y=115250
X512 11 VIA2_C_CDNS_7246542145924 $T=57320 145800 0 0 $X=57180 $Y=145090
X513 11 VIA2_C_CDNS_7246542145924 $T=58590 115960 0 0 $X=58450 $Y=115250
X514 11 VIA2_C_CDNS_7246542145924 $T=58590 145800 0 0 $X=58450 $Y=145090
X515 16 VIA2_C_CDNS_7246542145924 $T=59860 112400 0 0 $X=59720 $Y=111690
X516 17 VIA2_C_CDNS_7246542145924 $T=59860 149360 0 0 $X=59720 $Y=148650
X517 11 VIA2_C_CDNS_7246542145924 $T=60720 115960 0 0 $X=60580 $Y=115250
X518 11 VIA2_C_CDNS_7246542145924 $T=60720 145800 0 0 $X=60580 $Y=145090
X519 11 VIA2_C_CDNS_7246542145924 $T=61990 115960 0 0 $X=61850 $Y=115250
X520 11 VIA2_C_CDNS_7246542145924 $T=61990 145800 0 0 $X=61850 $Y=145090
X521 17 VIA2_C_CDNS_7246542145924 $T=63260 114180 0 0 $X=63120 $Y=113470
X522 16 VIA2_C_CDNS_7246542145924 $T=63260 147580 0 0 $X=63120 $Y=146870
X523 11 VIA2_C_CDNS_7246542145924 $T=64120 115960 0 0 $X=63980 $Y=115250
X524 11 VIA2_C_CDNS_7246542145924 $T=64120 145800 0 0 $X=63980 $Y=145090
X525 11 VIA2_C_CDNS_7246542145924 $T=65390 115960 0 0 $X=65250 $Y=115250
X526 11 VIA2_C_CDNS_7246542145924 $T=65390 145800 0 0 $X=65250 $Y=145090
X527 11 VIA2_C_CDNS_7246542145924 $T=66660 115960 0 0 $X=66520 $Y=115250
X528 11 VIA2_C_CDNS_7246542145924 $T=66660 145800 0 0 $X=66520 $Y=145090
X529 16 VIA3_C_CDNS_7246542145925 $T=7620 112400 0 0 $X=6910 $Y=111740
X530 16 VIA3_C_CDNS_7246542145925 $T=7620 147580 0 0 $X=6910 $Y=146920
X531 17 VIA3_C_CDNS_7246542145925 $T=9500 114180 0 0 $X=8790 $Y=113520
X532 17 VIA3_C_CDNS_7246542145925 $T=9500 149360 0 0 $X=8790 $Y=148700
X533 11 VIA3_C_CDNS_7246542145925 $T=11380 115960 0 0 $X=10670 $Y=115300
X534 11 VIA3_C_CDNS_7246542145925 $T=11380 145800 0 0 $X=10670 $Y=145140
X535 11 VIA3_C_CDNS_7246542145925 $T=68400 115960 0 0 $X=67690 $Y=115300
X536 11 VIA3_C_CDNS_7246542145925 $T=68400 145800 0 0 $X=67690 $Y=145140
X537 16 VIA3_C_CDNS_7246542145925 $T=70280 112400 0 0 $X=69570 $Y=111740
X538 16 VIA3_C_CDNS_7246542145925 $T=70280 147580 0 0 $X=69570 $Y=146920
X539 17 VIA3_C_CDNS_7246542145925 $T=72160 114180 0 0 $X=71450 $Y=113520
X540 17 VIA3_C_CDNS_7246542145925 $T=72160 149360 0 0 $X=71450 $Y=148700
X541 1 VIA1_C_CDNS_7246542145926 $T=15905 4500 0 0 $X=13335 $Y=3230
X542 1 VIA1_C_CDNS_7246542145926 $T=62500 4500 0 0 $X=59930 $Y=3230
X543 9 VIA2_C_CDNS_7246542145927 $T=17575 53125 0 0 $X=16825 $Y=52375
X544 13 VIA2_C_CDNS_7246542145927 $T=163125 148400 0 0 $X=162375 $Y=147650
X545 14 VIA2_C_CDNS_7246542145927 $T=204535 148400 0 0 $X=203785 $Y=147650
X546 15 VIA2_C_CDNS_7246542145927 $T=226740 148400 0 0 $X=225990 $Y=147650
X547 4 VIA2_C_CDNS_7246542145928 $T=170630 146620 0 0 $X=168580 $Y=145870
X548 6 VIA2_C_CDNS_7246542145928 $T=196715 146620 0 0 $X=194665 $Y=145870
X549 5 VIA2_C_CDNS_7246542145928 $T=220620 146620 0 0 $X=218570 $Y=145870
X550 18 VIA2_C_CDNS_7246542145936 $T=82800 119325 0 0 $X=82310 $Y=117275
X551 4 VIA2_C_CDNS_7246542145936 $T=82850 149150 0 0 $X=82360 $Y=147100
X552 18 VIA1_C_CDNS_7246542145937 $T=82800 119325 0 0 $X=82310 $Y=117275
X553 4 VIA1_C_CDNS_7246542145937 $T=82850 149150 0 0 $X=82360 $Y=147100
X554 2 1 VIA1_C_CDNS_7246542145940 $T=70935 208110 0 0 $X=65765 $Y=205540
X555 2 1 VIA1_C_CDNS_7246542145940 $T=150700 208200 0 0 $X=145530 $Y=205630
X556 14 8 6 2 1 pe3_CDNS_724654214590 $T=189280 150320 0 0 $X=187770 $Y=149290
X557 15 8 5 2 1 pe3_CDNS_724654214590 $T=213190 150320 0 0 $X=211680 $Y=149290
X558 1 1 1 ne3_CDNS_724654214591 $T=17980 14080 0 0 $X=17180 $Y=13680
X559 1 1 1 ne3_CDNS_724654214591 $T=17980 30170 0 0 $X=17180 $Y=29770
X560 1 9 10 ne3_CDNS_724654214591 $T=24220 14080 0 0 $X=23420 $Y=13680
X561 1 9 9 ne3_CDNS_724654214591 $T=24220 30170 0 0 $X=23420 $Y=29770
X562 1 9 9 ne3_CDNS_724654214591 $T=30460 14080 0 0 $X=29660 $Y=13680
X563 1 9 10 ne3_CDNS_724654214591 $T=30460 30170 0 0 $X=29660 $Y=29770
X564 1 9 8 ne3_CDNS_724654214591 $T=36700 14080 0 0 $X=35900 $Y=13680
X565 1 9 9 ne3_CDNS_724654214591 $T=36700 30170 0 0 $X=35900 $Y=29770
X566 1 9 9 ne3_CDNS_724654214591 $T=42940 14080 0 0 $X=42140 $Y=13680
X567 1 9 10 ne3_CDNS_724654214591 $T=42940 30170 0 0 $X=42140 $Y=29770
X568 1 9 10 ne3_CDNS_724654214591 $T=49180 14080 0 0 $X=48380 $Y=13680
X569 1 1 1 ne3_CDNS_724654214591 $T=49180 30170 0 0 $X=48380 $Y=29770
X570 1 1 1 ne3_CDNS_724654214591 $T=55420 14080 0 0 $X=54620 $Y=13680
X571 1 1 1 ne3_CDNS_724654214591 $T=55420 30170 0 0 $X=54620 $Y=29770
X572 13 8 4 2 1 pe3_CDNS_724654214592 $T=162340 150320 0 0 $X=160830 $Y=149290
X573 2 12 2 1 pe3_CDNS_724654214593 $T=138060 190125 0 0 $X=136550 $Y=189095
X574 12 8 2 1 pe3_CDNS_724654214593 $T=147620 190125 0 0 $X=146110 $Y=189095
X575 4 18 1 rpp1k1_3_CDNS_724654214594 $T=87870 117335 0 0 $X=82710 $Y=117115
X576 9 3 3 1 ne3_CDNS_724654214595 $T=17545 54415 0 0 $X=16745 $Y=54015
X577 10 3 11 1 ne3_CDNS_724654214595 $T=42480 54195 0 0 $X=41680 $Y=53795
X578 2 2 2 1 pe3_CDNS_724654214599 $T=165675 175935 0 0 $X=164165 $Y=174905
X579 2 2 2 1 pe3_CDNS_724654214599 $T=165675 195955 0 0 $X=164165 $Y=194925
X580 2 17 14 1 pe3_CDNS_724654214599 $T=168915 175935 0 0 $X=167405 $Y=174905
X581 2 17 15 1 pe3_CDNS_724654214599 $T=168915 195955 0 0 $X=167405 $Y=194925
X582 2 17 15 1 pe3_CDNS_724654214599 $T=172155 175935 0 0 $X=170645 $Y=174905
X583 2 17 13 1 pe3_CDNS_724654214599 $T=172155 195955 0 0 $X=170645 $Y=194925
X584 2 17 13 1 pe3_CDNS_724654214599 $T=175395 175935 0 0 $X=173885 $Y=174905
X585 2 17 14 1 pe3_CDNS_724654214599 $T=175395 195955 0 0 $X=173885 $Y=194925
X586 2 17 14 1 pe3_CDNS_724654214599 $T=178635 175935 0 0 $X=177125 $Y=174905
X587 2 17 15 1 pe3_CDNS_724654214599 $T=178635 195955 0 0 $X=177125 $Y=194925
X588 2 17 13 1 pe3_CDNS_724654214599 $T=181875 175935 0 0 $X=180365 $Y=174905
X589 2 17 15 1 pe3_CDNS_724654214599 $T=181875 195955 0 0 $X=180365 $Y=194925
X590 2 17 15 1 pe3_CDNS_724654214599 $T=185115 175935 0 0 $X=183605 $Y=174905
X591 2 17 13 1 pe3_CDNS_724654214599 $T=185115 195955 0 0 $X=183605 $Y=194925
X592 2 17 13 1 pe3_CDNS_724654214599 $T=188355 175935 0 0 $X=186845 $Y=174905
X593 2 17 14 1 pe3_CDNS_724654214599 $T=188355 195955 0 0 $X=186845 $Y=194925
X594 2 17 14 1 pe3_CDNS_724654214599 $T=191595 175935 0 0 $X=190085 $Y=174905
X595 2 17 13 1 pe3_CDNS_724654214599 $T=191595 195955 0 0 $X=190085 $Y=194925
X596 2 17 13 1 pe3_CDNS_724654214599 $T=194835 175935 0 0 $X=193325 $Y=174905
X597 2 17 15 1 pe3_CDNS_724654214599 $T=194835 195955 0 0 $X=193325 $Y=194925
X598 2 17 15 1 pe3_CDNS_724654214599 $T=198075 175935 0 0 $X=196565 $Y=174905
X599 2 17 13 1 pe3_CDNS_724654214599 $T=198075 195955 0 0 $X=196565 $Y=194925
X600 2 17 13 1 pe3_CDNS_724654214599 $T=201315 175935 0 0 $X=199805 $Y=174905
X601 2 17 14 1 pe3_CDNS_724654214599 $T=201315 195955 0 0 $X=199805 $Y=194925
X602 2 17 14 1 pe3_CDNS_724654214599 $T=204555 175935 0 0 $X=203045 $Y=174905
X603 2 17 13 1 pe3_CDNS_724654214599 $T=204555 195955 0 0 $X=203045 $Y=194925
X604 2 17 14 1 pe3_CDNS_724654214599 $T=207795 175935 0 0 $X=206285 $Y=174905
X605 2 17 15 1 pe3_CDNS_724654214599 $T=207795 195955 0 0 $X=206285 $Y=194925
X606 2 17 15 1 pe3_CDNS_724654214599 $T=211035 175935 0 0 $X=209525 $Y=174905
X607 2 17 13 1 pe3_CDNS_724654214599 $T=211035 195955 0 0 $X=209525 $Y=194925
X608 2 17 13 1 pe3_CDNS_724654214599 $T=214275 175935 0 0 $X=212765 $Y=174905
X609 2 17 14 1 pe3_CDNS_724654214599 $T=214275 195955 0 0 $X=212765 $Y=194925
X610 2 17 14 1 pe3_CDNS_724654214599 $T=217515 175935 0 0 $X=216005 $Y=174905
X611 2 17 15 1 pe3_CDNS_724654214599 $T=217515 195955 0 0 $X=216005 $Y=194925
X612 2 2 2 1 pe3_CDNS_724654214599 $T=220755 175935 0 0 $X=219245 $Y=174905
X613 2 2 2 1 pe3_CDNS_724654214599 $T=220755 195955 0 0 $X=219245 $Y=194925
X614 2 2 2 1 pe3_CDNS_7246542145910 $T=12010 172320 0 0 $X=10500 $Y=171290
X615 2 2 2 1 pe3_CDNS_7246542145910 $T=12010 190000 0 0 $X=10500 $Y=188970
X616 2 16 16 1 pe3_CDNS_7246542145910 $T=23250 172320 0 0 $X=21740 $Y=171290
X617 2 16 17 1 pe3_CDNS_7246542145910 $T=23250 190000 0 0 $X=21740 $Y=188970
X618 2 16 17 1 pe3_CDNS_7246542145910 $T=34490 172320 0 0 $X=32980 $Y=171290
X619 2 16 16 1 pe3_CDNS_7246542145910 $T=34490 190000 0 0 $X=32980 $Y=188970
X620 2 16 16 1 pe3_CDNS_7246542145910 $T=45730 172320 0 0 $X=44220 $Y=171290
X621 2 16 17 1 pe3_CDNS_7246542145910 $T=45730 190000 0 0 $X=44220 $Y=188970
X622 2 16 17 1 pe3_CDNS_7246542145910 $T=56970 172320 0 0 $X=55460 $Y=171290
X623 2 16 16 1 pe3_CDNS_7246542145910 $T=56970 190000 0 0 $X=55460 $Y=188970
X624 2 16 16 1 pe3_CDNS_7246542145910 $T=68210 172320 0 0 $X=66700 $Y=171290
X625 2 16 17 1 pe3_CDNS_7246542145910 $T=68210 190000 0 0 $X=66700 $Y=188970
X626 2 16 17 1 pe3_CDNS_7246542145910 $T=79450 172320 0 0 $X=77940 $Y=171290
X627 2 16 16 1 pe3_CDNS_7246542145910 $T=79450 190000 0 0 $X=77940 $Y=188970
X628 2 16 16 1 pe3_CDNS_7246542145910 $T=90690 172320 0 0 $X=89180 $Y=171290
X629 2 16 17 1 pe3_CDNS_7246542145910 $T=90690 190000 0 0 $X=89180 $Y=188970
X630 2 16 17 1 pe3_CDNS_7246542145910 $T=101930 172320 0 0 $X=100420 $Y=171290
X631 2 16 16 1 pe3_CDNS_7246542145910 $T=101930 190000 0 0 $X=100420 $Y=188970
X632 2 2 2 1 pe3_CDNS_7246542145910 $T=113170 172320 0 0 $X=111660 $Y=171290
X633 2 2 2 1 pe3_CDNS_7246542145910 $T=113170 190000 0 0 $X=111660 $Y=188970
X634 11 2 11 11 11 17 16 4 11 7
+ 1 MASCO__B5 $T=9330 114030 0 0 $X=9330 $Y=114030
X635 11 2 16 17 4 17 16 4 7 7
+ 1 MASCO__B5 $T=16130 114030 0 0 $X=16130 $Y=114030
X636 11 2 16 17 4 17 16 4 7 7
+ 1 MASCO__B5 $T=22930 114030 0 0 $X=22930 $Y=114030
X637 11 2 16 17 4 17 16 4 7 7
+ 1 MASCO__B5 $T=29730 114030 0 0 $X=29730 $Y=114030
X638 11 2 16 17 4 17 16 4 7 7
+ 1 MASCO__B5 $T=36530 114030 0 0 $X=36530 $Y=114030
X639 11 2 16 17 4 17 16 4 7 7
+ 1 MASCO__B5 $T=43330 114030 0 0 $X=43330 $Y=114030
X640 11 2 16 17 4 17 16 4 7 7
+ 1 MASCO__B5 $T=50130 114030 0 0 $X=50130 $Y=114030
X641 11 2 16 17 4 11 11 11 7 11
+ 1 MASCO__B5 $T=56930 114030 0 0 $X=56930 $Y=114030
X642 5 1 1 MOSVC3 w=3e-05 l=3e-05 $X=85530 $Y=8110 $dt=3
X643 5 1 1 MOSVC3 w=3e-05 l=3e-05 $X=85530 $Y=39350 $dt=3
X644 5 1 1 MOSVC3 w=3e-05 l=3e-05 $X=85530 $Y=70590 $dt=3
X645 6 1 1 MOSVC3 w=3e-05 l=3e-05 $X=122495 $Y=8050 $dt=3
X646 6 1 1 MOSVC3 w=3e-05 l=3e-05 $X=122495 $Y=39290 $dt=3
X647 6 1 1 MOSVC3 w=3e-05 l=3e-05 $X=122495 $Y=70530 $dt=3
D6 1 2 p_dnw AREA=2.36318e-09 PJ=0.00033402 perimeter=0.00033402 $X=4385 $Y=163650 $dt=5
D7 1 2 p_dnw AREA=2.57209e-10 PJ=8.388e-05 perimeter=8.388e-05 $X=134410 $Y=183535 $dt=5
D8 1 2 p_dnw AREA=1.81014e-09 PJ=0.00023539 perimeter=0.00023539 $X=158410 $Y=166295 $dt=5
D9 1 2 p_dnw AREA=8.15582e-10 PJ=0.0001871 perimeter=0.0001871 $X=158690 $Y=143730 $dt=5
D10 1 2 p_dnw AREA=9.45702e-09 PJ=0.00040696 perimeter=0.00040696 $X=159475 $Y=6005 $dt=5
D11 1 2 p_ddnw AREA=1.66704e-09 PJ=0.0001998 perimeter=0.0001998 $X=8060 $Y=112760 $dt=6
D12 11 2 p_dipdnwmv AREA=9.57098e-10 PJ=0.000169 perimeter=0.000169 $X=11910 $Y=116610 $dt=7
D13 1 2 p_dnw3 AREA=1.37701e-09 PJ=0 perimeter=0 $X=10500 $Y=171290 $dt=8
D14 1 2 p_dnw3 AREA=1.37701e-09 PJ=0 perimeter=0 $X=10500 $Y=188970 $dt=8
D15 1 1 p_dnw3 AREA=2.03309e-10 PJ=0.00024988 perimeter=0.00024988 $X=85100 $Y=7310 $dt=8
D16 1 1 p_dnw3 AREA=2.03309e-10 PJ=0.00024988 perimeter=0.00024988 $X=122065 $Y=7250 $dt=8
D17 1 2 p_dnw3 AREA=7.24806e-10 PJ=0 perimeter=0 $X=164165 $Y=174905 $dt=8
D18 1 2 p_dnw3 AREA=7.24806e-10 PJ=0 perimeter=0 $X=164165 $Y=194925 $dt=8
C19 17 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=161615 $Y=8145 $dt=11
C20 17 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=161615 $Y=39745 $dt=11
C21 17 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=161615 $Y=71345 $dt=11
C22 17 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=161615 $Y=102945 $dt=11
C23 17 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=196615 $Y=8145 $dt=11
C24 17 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=196615 $Y=39745 $dt=11
C25 17 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=196615 $Y=71345 $dt=11
C26 17 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=196615 $Y=102945 $dt=11
.ends ref_bias

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246542145944                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246542145944 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246542145944

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246542145946                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246542145946 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246542145946

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246542145947                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246542145947 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246542145947

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246542145949                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246542145949 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246542145949

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246542145951                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246542145951 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246542145951

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246542145957                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246542145957 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246542145957

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246542145958                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246542145958 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246542145958

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246542145959                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246542145959 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246542145959

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246542145911                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246542145911 1 2 3 4 5
** N=5 EP=5 FDC=5
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=1
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=1
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=1
D4 5 4 p_dnw3 AREA=1.04198e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=8
.ends pe3_CDNS_7246542145911

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7246542145912                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7246542145912 1 2 3 4
** N=4 EP=4 FDC=4
M0 3 2 1 4 ne3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
M1 1 2 3 4 ne3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=0
M2 3 2 1 4 ne3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=0
M3 1 2 3 4 ne3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=0
.ends ne3_CDNS_7246542145912

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7246542145913                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7246542145913 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.0005215 W=8e-06 $[rpp1k1_3] $SUB=3 $X=-8220 $Y=0 $dt=9
.ends rpp1k1_3_CDNS_7246542145913

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7246542145914                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7246542145914 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.00082283 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=9
.ends rpp1k1_3_CDNS_7246542145914

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7246542145915                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7246542145915 1 2 3 4
** N=4 EP=4 FDC=1
M0 3 2 1 4 ne3 L=1e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
.ends ne3_CDNS_7246542145915

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246542145916                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246542145916 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=1
M0 3 2 1 4 pe3 L=5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_7246542145916

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246542145917                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246542145917 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 3 2 1 4 pe3 L=5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
D1 5 4 p_dnw3 AREA=9.67212e-11 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=8
.ends pe3_CDNS_7246542145917

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7246542145918                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7246542145918 1 2 3
** N=3 EP=3 FDC=1
M0 2 2 1 3 ne3 L=2e-06 W=1e-06 AD=4.8e-13 AS=4.8e-13 PD=2.96e-06 PS=2.96e-06 $X=0 $Y=0 $dt=0
.ends ne3_CDNS_7246542145918

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246542145919                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246542145919 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
M0 3 2 1 1 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_7246542145919

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7246542145920                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7246542145920 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.00082283 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=9
.ends rpp1k1_3_CDNS_7246542145920

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: bandgap_su                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt bandgap_su 1 2 3 4
** N=24 EP=4 FDC=165
X0 5 VIA2_C_CDNS_724654214590 $T=26170 76265 0 0 $X=25420 $Y=75515
X1 6 VIA1_C_CDNS_724654214597 $T=10135 89745 0 0 $X=9995 $Y=89555
X2 3 VIA1_C_CDNS_724654214597 $T=10845 66505 0 0 $X=10705 $Y=66315
X3 6 VIA1_C_CDNS_724654214597 $T=11675 89745 0 0 $X=11535 $Y=89555
X4 3 VIA1_C_CDNS_724654214597 $T=12385 66505 0 0 $X=12245 $Y=66315
X5 6 VIA1_C_CDNS_724654214597 $T=13215 89745 0 0 $X=13075 $Y=89555
X6 3 VIA1_C_CDNS_724654214597 $T=13925 66505 0 0 $X=13785 $Y=66315
X7 6 VIA1_C_CDNS_724654214597 $T=14755 89745 0 0 $X=14615 $Y=89555
X8 3 VIA1_C_CDNS_724654214597 $T=15465 66505 0 0 $X=15325 $Y=66315
X9 7 VIA1_C_CDNS_724654214597 $T=15870 27855 0 0 $X=15730 $Y=27665
X10 7 VIA1_C_CDNS_724654214597 $T=18110 27855 0 0 $X=17970 $Y=27665
X11 7 VIA1_C_CDNS_724654214597 $T=20350 27855 0 0 $X=20210 $Y=27665
X12 7 VIA1_C_CDNS_724654214597 $T=22590 27855 0 0 $X=22450 $Y=27665
X13 3 VIA1_C_CDNS_724654214597 $T=23230 66505 0 0 $X=23090 $Y=66315
X14 3 VIA1_C_CDNS_724654214597 $T=24770 66505 0 0 $X=24630 $Y=66315
X15 7 VIA1_C_CDNS_724654214597 $T=24830 27855 0 0 $X=24690 $Y=27665
X16 3 VIA1_C_CDNS_724654214597 $T=26310 66505 0 0 $X=26170 $Y=66315
X17 3 VIA1_C_CDNS_724654214597 $T=27850 66505 0 0 $X=27710 $Y=66315
X18 8 VIA1_C_CDNS_724654214599 $T=13400 117700 0 0 $X=13000 $Y=117510
X19 8 VIA1_C_CDNS_724654214599 $T=15640 117700 0 0 $X=15240 $Y=117510
X20 8 VIA1_C_CDNS_724654214599 $T=17880 117700 0 0 $X=17480 $Y=117510
X21 8 VIA1_C_CDNS_724654214599 $T=20120 117700 0 0 $X=19720 $Y=117510
X22 8 VIA1_C_CDNS_724654214599 $T=22360 117700 0 0 $X=21960 $Y=117510
X23 6 VIA1_C_CDNS_724654214599 $T=23940 89745 0 0 $X=23540 $Y=89555
X24 8 VIA1_C_CDNS_724654214599 $T=24600 117700 0 0 $X=24200 $Y=117510
X25 6 VIA1_C_CDNS_724654214599 $T=25480 89745 0 0 $X=25080 $Y=89555
X26 8 VIA1_C_CDNS_724654214599 $T=26840 117700 0 0 $X=26440 $Y=117510
X27 6 VIA1_C_CDNS_724654214599 $T=27020 89745 0 0 $X=26620 $Y=89555
X28 6 VIA1_C_CDNS_724654214599 $T=28560 89745 0 0 $X=28160 $Y=89555
X29 8 VIA1_C_CDNS_724654214599 $T=29080 117700 0 0 $X=28680 $Y=117510
X30 8 VIA1_C_CDNS_724654214599 $T=31320 117700 0 0 $X=30920 $Y=117510
X31 8 VIA1_C_CDNS_724654214599 $T=33560 117700 0 0 $X=33160 $Y=117510
X32 8 VIA1_C_CDNS_724654214599 $T=35800 117700 0 0 $X=35400 $Y=117510
X33 8 VIA1_C_CDNS_724654214599 $T=38040 117700 0 0 $X=37640 $Y=117510
X34 9 VIA1_C_CDNS_724654214599 $T=51305 71565 0 0 $X=50905 $Y=71375
X35 10 VIA1_C_CDNS_724654214599 $T=52955 72345 0 0 $X=52555 $Y=72155
X36 11 VIA1_C_CDNS_724654214599 $T=53520 26400 0 0 $X=53120 $Y=26210
X37 9 VIA1_C_CDNS_724654214599 $T=58085 71565 0 0 $X=57685 $Y=71375
X38 10 VIA1_C_CDNS_724654214599 $T=58765 72345 0 0 $X=58365 $Y=72155
X39 11 VIA1_C_CDNS_724654214599 $T=59760 26400 0 0 $X=59360 $Y=26210
X40 12 VIA1_C_CDNS_724654214599 $T=62155 117840 0 0 $X=61755 $Y=117650
X41 9 VIA1_C_CDNS_724654214599 $T=63785 71565 0 0 $X=63385 $Y=71375
X42 10 VIA1_C_CDNS_724654214599 $T=65435 72345 0 0 $X=65035 $Y=72155
X43 11 VIA1_C_CDNS_724654214599 $T=66000 26400 0 0 $X=65600 $Y=26210
X44 12 VIA1_C_CDNS_724654214599 $T=68395 117840 0 0 $X=67995 $Y=117650
X45 9 VIA1_C_CDNS_724654214599 $T=70565 71565 0 0 $X=70165 $Y=71375
X46 10 VIA1_C_CDNS_724654214599 $T=71245 72345 0 0 $X=70845 $Y=72155
X47 11 VIA1_C_CDNS_724654214599 $T=72240 26400 0 0 $X=71840 $Y=26210
X48 9 VIA1_C_CDNS_724654214599 $T=76265 71565 0 0 $X=75865 $Y=71375
X49 10 VIA1_C_CDNS_724654214599 $T=77915 72345 0 0 $X=77515 $Y=72155
X50 11 VIA1_C_CDNS_724654214599 $T=78480 26400 0 0 $X=78080 $Y=26210
X51 13 VIA1_C_CDNS_724654214599 $T=81575 136880 0 0 $X=81175 $Y=136690
X52 9 VIA1_C_CDNS_724654214599 $T=83045 71565 0 0 $X=82645 $Y=71375
X53 10 VIA1_C_CDNS_724654214599 $T=83725 72345 0 0 $X=83325 $Y=72155
X54 11 VIA1_C_CDNS_724654214599 $T=84720 26400 0 0 $X=84320 $Y=26210
X55 13 VIA1_C_CDNS_724654214599 $T=87815 136880 0 0 $X=87415 $Y=136690
X56 9 VIA1_C_CDNS_724654214599 $T=88745 71565 0 0 $X=88345 $Y=71375
X57 10 VIA1_C_CDNS_724654214599 $T=90395 72345 0 0 $X=89995 $Y=72155
X58 11 VIA1_C_CDNS_724654214599 $T=90960 26400 0 0 $X=90560 $Y=26210
X59 9 VIA1_C_CDNS_724654214599 $T=95525 71565 0 0 $X=95125 $Y=71375
X60 10 VIA1_C_CDNS_724654214599 $T=96205 72345 0 0 $X=95805 $Y=72155
X61 14 VIA1_C_CDNS_724654214599 $T=96290 114275 0 0 $X=95890 $Y=114085
X62 11 VIA1_C_CDNS_724654214599 $T=97200 26400 0 0 $X=96800 $Y=26210
X63 14 VIA1_C_CDNS_724654214599 $T=97830 114275 0 0 $X=97430 $Y=114085
X64 4 VIA1_C_CDNS_724654214599 $T=98460 136920 0 0 $X=98060 $Y=136730
X65 14 VIA1_C_CDNS_724654214599 $T=99370 114275 0 0 $X=98970 $Y=114085
X66 15 VIA1_C_CDNS_724654214599 $T=100700 136140 0 0 $X=100300 $Y=135950
X67 14 VIA1_C_CDNS_724654214599 $T=100910 114275 0 0 $X=100510 $Y=114085
X68 8 VIA1_C_CDNS_7246542145912 $T=9365 74485 0 0 $X=9225 $Y=73775
X69 7 VIA1_C_CDNS_7246542145912 $T=10075 52335 0 0 $X=9935 $Y=51625
X70 2 VIA1_C_CDNS_7246542145912 $T=10390 104220 0 0 $X=10250 $Y=103510
X71 2 VIA1_C_CDNS_7246542145912 $T=10390 131040 0 0 $X=10250 $Y=130330
X72 6 VIA1_C_CDNS_7246542145912 $T=10905 76265 0 0 $X=10765 $Y=75555
X73 3 VIA1_C_CDNS_7246542145912 $T=11615 54115 0 0 $X=11475 $Y=53405
X74 2 VIA1_C_CDNS_7246542145912 $T=11930 104220 0 0 $X=11790 $Y=103510
X75 2 VIA1_C_CDNS_7246542145912 $T=11930 131040 0 0 $X=11790 $Y=130330
X76 8 VIA1_C_CDNS_7246542145912 $T=12445 74485 0 0 $X=12305 $Y=73775
X77 2 VIA1_C_CDNS_7246542145912 $T=12630 104220 0 0 $X=12490 $Y=103510
X78 2 VIA1_C_CDNS_7246542145912 $T=12630 131040 0 0 $X=12490 $Y=130330
X79 1 VIA1_C_CDNS_7246542145912 $T=12860 15465 0 0 $X=12720 $Y=14755
X80 1 VIA1_C_CDNS_7246542145912 $T=12860 40105 0 0 $X=12720 $Y=39395
X81 7 VIA1_C_CDNS_7246542145912 $T=13155 52335 0 0 $X=13015 $Y=51625
X82 6 VIA1_C_CDNS_7246542145912 $T=13985 76265 0 0 $X=13845 $Y=75555
X83 4 VIA1_C_CDNS_7246542145912 $T=14170 98880 0 0 $X=14030 $Y=98170
X84 4 VIA1_C_CDNS_7246542145912 $T=14170 132820 0 0 $X=14030 $Y=132110
X85 1 VIA1_C_CDNS_7246542145912 $T=14400 15465 0 0 $X=14260 $Y=14755
X86 1 VIA1_C_CDNS_7246542145912 $T=14400 40105 0 0 $X=14260 $Y=39395
X87 3 VIA1_C_CDNS_7246542145912 $T=14695 54115 0 0 $X=14555 $Y=53405
X88 2 VIA1_C_CDNS_7246542145912 $T=14870 104220 0 0 $X=14730 $Y=103510
X89 2 VIA1_C_CDNS_7246542145912 $T=14870 131040 0 0 $X=14730 $Y=130330
X90 1 VIA1_C_CDNS_7246542145912 $T=15100 15465 0 0 $X=14960 $Y=14755
X91 1 VIA1_C_CDNS_7246542145912 $T=15100 40105 0 0 $X=14960 $Y=39395
X92 8 VIA1_C_CDNS_7246542145912 $T=15525 74485 0 0 $X=15385 $Y=73775
X93 7 VIA1_C_CDNS_7246542145912 $T=16235 52335 0 0 $X=16095 $Y=51625
X94 4 VIA1_C_CDNS_7246542145912 $T=16410 98880 0 0 $X=16270 $Y=98170
X95 4 VIA1_C_CDNS_7246542145912 $T=16410 132820 0 0 $X=16270 $Y=132110
X96 16 VIA1_C_CDNS_7246542145912 $T=16640 11905 0 0 $X=16500 $Y=11195
X97 7 VIA1_C_CDNS_7246542145912 $T=16640 43665 0 0 $X=16500 $Y=42955
X98 2 VIA1_C_CDNS_7246542145912 $T=17110 104220 0 0 $X=16970 $Y=103510
X99 2 VIA1_C_CDNS_7246542145912 $T=17110 131040 0 0 $X=16970 $Y=130330
X100 1 VIA1_C_CDNS_7246542145912 $T=17340 15465 0 0 $X=17200 $Y=14755
X101 1 VIA1_C_CDNS_7246542145912 $T=17340 40105 0 0 $X=17200 $Y=39395
X102 5 VIA1_C_CDNS_7246542145912 $T=18650 102440 0 0 $X=18510 $Y=101730
X103 8 VIA1_C_CDNS_7246542145912 $T=18650 134600 0 0 $X=18510 $Y=133890
X104 7 VIA1_C_CDNS_7246542145912 $T=18880 13685 0 0 $X=18740 $Y=12975
X105 16 VIA1_C_CDNS_7246542145912 $T=18880 41885 0 0 $X=18740 $Y=41175
X106 2 VIA1_C_CDNS_7246542145912 $T=19350 104220 0 0 $X=19210 $Y=103510
X107 2 VIA1_C_CDNS_7246542145912 $T=19350 131040 0 0 $X=19210 $Y=130330
X108 1 VIA1_C_CDNS_7246542145912 $T=19580 15465 0 0 $X=19440 $Y=14755
X109 1 VIA1_C_CDNS_7246542145912 $T=19580 40105 0 0 $X=19440 $Y=39395
X110 4 VIA1_C_CDNS_7246542145912 $T=20890 98880 0 0 $X=20750 $Y=98170
X111 4 VIA1_C_CDNS_7246542145912 $T=20890 132820 0 0 $X=20750 $Y=132110
X112 17 VIA1_C_CDNS_7246542145912 $T=21120 10125 0 0 $X=20980 $Y=9415
X113 18 VIA1_C_CDNS_7246542145912 $T=21120 45445 0 0 $X=20980 $Y=44735
X114 2 VIA1_C_CDNS_7246542145912 $T=21590 104220 0 0 $X=21450 $Y=103510
X115 2 VIA1_C_CDNS_7246542145912 $T=21590 131040 0 0 $X=21450 $Y=130330
X116 1 VIA1_C_CDNS_7246542145912 $T=21820 15465 0 0 $X=21680 $Y=14755
X117 1 VIA1_C_CDNS_7246542145912 $T=21820 40105 0 0 $X=21680 $Y=39395
X118 16 VIA1_C_CDNS_7246542145912 $T=22460 54255 0 0 $X=22320 $Y=53545
X119 4 VIA1_C_CDNS_7246542145912 $T=23130 98880 0 0 $X=22990 $Y=98170
X120 4 VIA1_C_CDNS_7246542145912 $T=23130 132820 0 0 $X=22990 $Y=132110
X121 5 VIA1_C_CDNS_7246542145912 $T=23170 76265 0 0 $X=23030 $Y=75555
X122 16 VIA1_C_CDNS_7246542145912 $T=23360 11905 0 0 $X=23220 $Y=11195
X123 7 VIA1_C_CDNS_7246542145912 $T=23360 43665 0 0 $X=23220 $Y=42955
X124 2 VIA1_C_CDNS_7246542145912 $T=23830 104220 0 0 $X=23690 $Y=103510
X125 2 VIA1_C_CDNS_7246542145912 $T=23830 131040 0 0 $X=23690 $Y=130330
X126 6 VIA1_C_CDNS_7246542145912 $T=24000 52475 0 0 $X=23860 $Y=51765
X127 1 VIA1_C_CDNS_7246542145912 $T=24060 15465 0 0 $X=23920 $Y=14755
X128 1 VIA1_C_CDNS_7246542145912 $T=24060 40105 0 0 $X=23920 $Y=39395
X129 19 VIA1_C_CDNS_7246542145912 $T=24710 74485 0 0 $X=24570 $Y=73775
X130 8 VIA1_C_CDNS_7246542145912 $T=25370 100660 0 0 $X=25230 $Y=99950
X131 5 VIA1_C_CDNS_7246542145912 $T=25370 136380 0 0 $X=25230 $Y=135670
X132 16 VIA1_C_CDNS_7246542145912 $T=25540 54255 0 0 $X=25400 $Y=53545
X133 7 VIA1_C_CDNS_7246542145912 $T=25600 13685 0 0 $X=25460 $Y=12975
X134 16 VIA1_C_CDNS_7246542145912 $T=25600 41885 0 0 $X=25460 $Y=41175
X135 2 VIA1_C_CDNS_7246542145912 $T=26070 104220 0 0 $X=25930 $Y=103510
X136 2 VIA1_C_CDNS_7246542145912 $T=26070 131040 0 0 $X=25930 $Y=130330
X137 5 VIA1_C_CDNS_7246542145912 $T=26250 76265 0 0 $X=26110 $Y=75555
X138 1 VIA1_C_CDNS_7246542145912 $T=26300 15465 0 0 $X=26160 $Y=14755
X139 1 VIA1_C_CDNS_7246542145912 $T=26300 40105 0 0 $X=26160 $Y=39395
X140 6 VIA1_C_CDNS_7246542145912 $T=27080 52475 0 0 $X=26940 $Y=51765
X141 5 VIA1_C_CDNS_7246542145912 $T=27610 102440 0 0 $X=27470 $Y=101730
X142 8 VIA1_C_CDNS_7246542145912 $T=27610 134600 0 0 $X=27470 $Y=133890
X143 19 VIA1_C_CDNS_7246542145912 $T=27790 74485 0 0 $X=27650 $Y=73775
X144 1 VIA1_C_CDNS_7246542145912 $T=27840 15465 0 0 $X=27700 $Y=14755
X145 1 VIA1_C_CDNS_7246542145912 $T=27840 40105 0 0 $X=27700 $Y=39395
X146 2 VIA1_C_CDNS_7246542145912 $T=28310 104220 0 0 $X=28170 $Y=103510
X147 2 VIA1_C_CDNS_7246542145912 $T=28310 131040 0 0 $X=28170 $Y=130330
X148 16 VIA1_C_CDNS_7246542145912 $T=28620 54255 0 0 $X=28480 $Y=53545
X149 5 VIA1_C_CDNS_7246542145912 $T=29330 76265 0 0 $X=29190 $Y=75555
X150 4 VIA1_C_CDNS_7246542145912 $T=29850 98880 0 0 $X=29710 $Y=98170
X151 4 VIA1_C_CDNS_7246542145912 $T=29850 132820 0 0 $X=29710 $Y=132110
X152 2 VIA1_C_CDNS_7246542145912 $T=30550 104220 0 0 $X=30410 $Y=103510
X153 2 VIA1_C_CDNS_7246542145912 $T=30550 131040 0 0 $X=30410 $Y=130330
X154 4 VIA1_C_CDNS_7246542145912 $T=32090 98880 0 0 $X=31950 $Y=98170
X155 4 VIA1_C_CDNS_7246542145912 $T=32090 132820 0 0 $X=31950 $Y=132110
X156 2 VIA1_C_CDNS_7246542145912 $T=32790 104220 0 0 $X=32650 $Y=103510
X157 2 VIA1_C_CDNS_7246542145912 $T=32790 131040 0 0 $X=32650 $Y=130330
X158 8 VIA1_C_CDNS_7246542145912 $T=34330 100660 0 0 $X=34190 $Y=99950
X159 5 VIA1_C_CDNS_7246542145912 $T=34330 136380 0 0 $X=34190 $Y=135670
X160 2 VIA1_C_CDNS_7246542145912 $T=35030 104220 0 0 $X=34890 $Y=103510
X161 2 VIA1_C_CDNS_7246542145912 $T=35030 131040 0 0 $X=34890 $Y=130330
X162 4 VIA1_C_CDNS_7246542145912 $T=36570 98880 0 0 $X=36430 $Y=98170
X163 4 VIA1_C_CDNS_7246542145912 $T=36570 132820 0 0 $X=36430 $Y=132110
X164 2 VIA1_C_CDNS_7246542145912 $T=37270 104220 0 0 $X=37130 $Y=103510
X165 2 VIA1_C_CDNS_7246542145912 $T=37270 131040 0 0 $X=37130 $Y=130330
X166 4 VIA1_C_CDNS_7246542145912 $T=38810 98880 0 0 $X=38670 $Y=98170
X167 4 VIA1_C_CDNS_7246542145912 $T=38810 132820 0 0 $X=38670 $Y=132110
X168 2 VIA1_C_CDNS_7246542145912 $T=39510 104220 0 0 $X=39370 $Y=103510
X169 2 VIA1_C_CDNS_7246542145912 $T=39510 131040 0 0 $X=39370 $Y=130330
X170 2 VIA1_C_CDNS_7246542145912 $T=41050 104220 0 0 $X=40910 $Y=103510
X171 2 VIA1_C_CDNS_7246542145912 $T=41050 131040 0 0 $X=40910 $Y=130330
X172 19 VIA1_C_CDNS_7246542145912 $T=42835 58225 0 0 $X=42695 $Y=57515
X173 19 VIA1_C_CDNS_7246542145912 $T=42835 85685 0 0 $X=42695 $Y=84975
X174 1 VIA1_C_CDNS_7246542145912 $T=44510 14010 0 0 $X=44370 $Y=13300
X175 1 VIA1_C_CDNS_7246542145912 $T=44510 38730 0 0 $X=44370 $Y=38020
X176 19 VIA1_C_CDNS_7246542145912 $T=48375 58225 0 0 $X=48235 $Y=57515
X177 19 VIA1_C_CDNS_7246542145912 $T=48375 85685 0 0 $X=48235 $Y=84975
X178 19 VIA1_C_CDNS_7246542145912 $T=49075 58225 0 0 $X=48935 $Y=57515
X179 19 VIA1_C_CDNS_7246542145912 $T=49075 85685 0 0 $X=48935 $Y=84975
X180 1 VIA1_C_CDNS_7246542145912 $T=50050 14010 0 0 $X=49910 $Y=13300
X181 1 VIA1_C_CDNS_7246542145912 $T=50050 38730 0 0 $X=49910 $Y=38020
X182 1 VIA1_C_CDNS_7246542145912 $T=50750 14010 0 0 $X=50610 $Y=13300
X183 1 VIA1_C_CDNS_7246542145912 $T=50750 38730 0 0 $X=50610 $Y=38020
X184 14 VIA1_C_CDNS_7246542145912 $T=54615 54665 0 0 $X=54475 $Y=53955
X185 11 VIA1_C_CDNS_7246542145912 $T=54615 89245 0 0 $X=54475 $Y=88535
X186 19 VIA1_C_CDNS_7246542145912 $T=55315 58225 0 0 $X=55175 $Y=57515
X187 19 VIA1_C_CDNS_7246542145912 $T=55315 85685 0 0 $X=55175 $Y=84975
X188 11 VIA1_C_CDNS_7246542145912 $T=56290 12230 0 0 $X=56150 $Y=11520
X189 14 VIA1_C_CDNS_7246542145912 $T=56290 40510 0 0 $X=56150 $Y=39800
X190 1 VIA1_C_CDNS_7246542145912 $T=56990 14010 0 0 $X=56850 $Y=13300
X191 1 VIA1_C_CDNS_7246542145912 $T=56990 38730 0 0 $X=56850 $Y=38020
X192 11 VIA1_C_CDNS_7246542145912 $T=60855 56445 0 0 $X=60715 $Y=55735
X193 14 VIA1_C_CDNS_7246542145912 $T=60855 87465 0 0 $X=60715 $Y=86755
X194 19 VIA1_C_CDNS_7246542145912 $T=61555 58225 0 0 $X=61415 $Y=57515
X195 19 VIA1_C_CDNS_7246542145912 $T=61555 85685 0 0 $X=61415 $Y=84975
X196 14 VIA1_C_CDNS_7246542145912 $T=62530 10450 0 0 $X=62390 $Y=9740
X197 11 VIA1_C_CDNS_7246542145912 $T=62530 42290 0 0 $X=62390 $Y=41580
X198 1 VIA1_C_CDNS_7246542145912 $T=63230 14010 0 0 $X=63090 $Y=13300
X199 1 VIA1_C_CDNS_7246542145912 $T=63230 38730 0 0 $X=63090 $Y=38020
X200 14 VIA1_C_CDNS_7246542145912 $T=67095 54665 0 0 $X=66955 $Y=53955
X201 11 VIA1_C_CDNS_7246542145912 $T=67095 89245 0 0 $X=66955 $Y=88535
X202 19 VIA1_C_CDNS_7246542145912 $T=67795 58225 0 0 $X=67655 $Y=57515
X203 19 VIA1_C_CDNS_7246542145912 $T=67795 85685 0 0 $X=67655 $Y=84975
X204 11 VIA1_C_CDNS_7246542145912 $T=68770 12230 0 0 $X=68630 $Y=11520
X205 14 VIA1_C_CDNS_7246542145912 $T=68770 40510 0 0 $X=68630 $Y=39800
X206 1 VIA1_C_CDNS_7246542145912 $T=69470 14010 0 0 $X=69330 $Y=13300
X207 1 VIA1_C_CDNS_7246542145912 $T=69470 38730 0 0 $X=69330 $Y=38020
X208 11 VIA1_C_CDNS_7246542145912 $T=73335 56445 0 0 $X=73195 $Y=55735
X209 14 VIA1_C_CDNS_7246542145912 $T=73335 87465 0 0 $X=73195 $Y=86755
X210 19 VIA1_C_CDNS_7246542145912 $T=74035 58225 0 0 $X=73895 $Y=57515
X211 19 VIA1_C_CDNS_7246542145912 $T=74035 85685 0 0 $X=73895 $Y=84975
X212 14 VIA1_C_CDNS_7246542145912 $T=75010 10450 0 0 $X=74870 $Y=9740
X213 11 VIA1_C_CDNS_7246542145912 $T=75010 42290 0 0 $X=74870 $Y=41580
X214 1 VIA1_C_CDNS_7246542145912 $T=75710 14010 0 0 $X=75570 $Y=13300
X215 1 VIA1_C_CDNS_7246542145912 $T=75710 38730 0 0 $X=75570 $Y=38020
X216 2 VIA1_C_CDNS_7246542145912 $T=78805 123400 0 0 $X=78665 $Y=122690
X217 14 VIA1_C_CDNS_7246542145912 $T=79575 54665 0 0 $X=79435 $Y=53955
X218 11 VIA1_C_CDNS_7246542145912 $T=79575 89245 0 0 $X=79435 $Y=88535
X219 19 VIA1_C_CDNS_7246542145912 $T=80275 58225 0 0 $X=80135 $Y=57515
X220 19 VIA1_C_CDNS_7246542145912 $T=80275 85685 0 0 $X=80135 $Y=84975
X221 11 VIA1_C_CDNS_7246542145912 $T=81250 12230 0 0 $X=81110 $Y=11520
X222 14 VIA1_C_CDNS_7246542145912 $T=81250 40510 0 0 $X=81110 $Y=39800
X223 1 VIA1_C_CDNS_7246542145912 $T=81950 14010 0 0 $X=81810 $Y=13300
X224 1 VIA1_C_CDNS_7246542145912 $T=81950 38730 0 0 $X=81810 $Y=38020
X225 13 VIA1_C_CDNS_7246542145912 $T=84345 121620 0 0 $X=84205 $Y=120910
X226 2 VIA1_C_CDNS_7246542145912 $T=85045 123400 0 0 $X=84905 $Y=122690
X227 11 VIA1_C_CDNS_7246542145912 $T=85815 56445 0 0 $X=85675 $Y=55735
X228 14 VIA1_C_CDNS_7246542145912 $T=85815 87465 0 0 $X=85675 $Y=86755
X229 19 VIA1_C_CDNS_7246542145912 $T=86515 58225 0 0 $X=86375 $Y=57515
X230 19 VIA1_C_CDNS_7246542145912 $T=86515 85685 0 0 $X=86375 $Y=84975
X231 14 VIA1_C_CDNS_7246542145912 $T=87490 10450 0 0 $X=87350 $Y=9740
X232 11 VIA1_C_CDNS_7246542145912 $T=87490 42290 0 0 $X=87350 $Y=41580
X233 1 VIA1_C_CDNS_7246542145912 $T=88190 14010 0 0 $X=88050 $Y=13300
X234 1 VIA1_C_CDNS_7246542145912 $T=88190 38730 0 0 $X=88050 $Y=38020
X235 20 VIA1_C_CDNS_7246542145912 $T=90585 119840 0 0 $X=90445 $Y=119130
X236 14 VIA1_C_CDNS_7246542145912 $T=92055 54665 0 0 $X=91915 $Y=53955
X237 11 VIA1_C_CDNS_7246542145912 $T=92055 89245 0 0 $X=91915 $Y=88535
X238 19 VIA1_C_CDNS_7246542145912 $T=92755 58225 0 0 $X=92615 $Y=57515
X239 19 VIA1_C_CDNS_7246542145912 $T=92755 85685 0 0 $X=92615 $Y=84975
X240 11 VIA1_C_CDNS_7246542145912 $T=93730 12230 0 0 $X=93590 $Y=11520
X241 14 VIA1_C_CDNS_7246542145912 $T=93730 40510 0 0 $X=93590 $Y=39800
X242 1 VIA1_C_CDNS_7246542145912 $T=94430 14010 0 0 $X=94290 $Y=13300
X243 1 VIA1_C_CDNS_7246542145912 $T=94430 38730 0 0 $X=94290 $Y=38020
X244 11 VIA1_C_CDNS_7246542145912 $T=98295 56445 0 0 $X=98155 $Y=55735
X245 14 VIA1_C_CDNS_7246542145912 $T=98295 87465 0 0 $X=98155 $Y=86755
X246 19 VIA1_C_CDNS_7246542145912 $T=98995 58225 0 0 $X=98855 $Y=57515
X247 19 VIA1_C_CDNS_7246542145912 $T=98995 85685 0 0 $X=98855 $Y=84975
X248 14 VIA1_C_CDNS_7246542145912 $T=99970 10450 0 0 $X=99830 $Y=9740
X249 11 VIA1_C_CDNS_7246542145912 $T=99970 42290 0 0 $X=99830 $Y=41580
X250 1 VIA1_C_CDNS_7246542145912 $T=100670 14010 0 0 $X=100530 $Y=13300
X251 1 VIA1_C_CDNS_7246542145912 $T=100670 38730 0 0 $X=100530 $Y=38020
X252 19 VIA1_C_CDNS_7246542145912 $T=104535 58225 0 0 $X=104395 $Y=57515
X253 19 VIA1_C_CDNS_7246542145912 $T=104535 85685 0 0 $X=104395 $Y=84975
X254 1 VIA1_C_CDNS_7246542145912 $T=106210 14010 0 0 $X=106070 $Y=13300
X255 1 VIA1_C_CDNS_7246542145912 $T=106210 38730 0 0 $X=106070 $Y=38020
X256 8 VIA2_C_CDNS_7246542145913 $T=5840 117700 0 0 $X=5130 $Y=117560
X257 7 VIA2_C_CDNS_7246542145913 $T=7240 27855 0 0 $X=6530 $Y=27715
X258 2 VIA2_C_CDNS_7246542145918 $T=7870 104220 0 0 $X=6900 $Y=103560
X259 2 VIA2_C_CDNS_7246542145918 $T=7870 131040 0 0 $X=6900 $Y=130380
X260 1 VIA2_C_CDNS_7246542145918 $T=11050 15465 0 0 $X=10080 $Y=14805
X261 1 VIA2_C_CDNS_7246542145918 $T=11050 40105 0 0 $X=10080 $Y=39445
X262 1 VIA2_C_CDNS_7246542145918 $T=29650 15465 0 0 $X=28680 $Y=14805
X263 1 VIA2_C_CDNS_7246542145918 $T=29650 40105 0 0 $X=28680 $Y=39445
X264 11 VIA2_C_CDNS_7246542145918 $T=38035 56445 0 0 $X=37065 $Y=55785
X265 11 VIA2_C_CDNS_7246542145918 $T=38035 89245 0 0 $X=37065 $Y=88585
X266 19 VIA2_C_CDNS_7246542145918 $T=40315 58225 0 0 $X=39345 $Y=57565
X267 19 VIA2_C_CDNS_7246542145918 $T=40315 85685 0 0 $X=39345 $Y=85025
X268 11 VIA2_C_CDNS_7246542145918 $T=40420 12230 0 0 $X=39450 $Y=11570
X269 11 VIA2_C_CDNS_7246542145918 $T=40420 42290 0 0 $X=39450 $Y=41630
X270 1 VIA2_C_CDNS_7246542145918 $T=42700 14010 0 0 $X=41730 $Y=13350
X271 1 VIA2_C_CDNS_7246542145918 $T=42700 38730 0 0 $X=41730 $Y=38070
X272 2 VIA2_C_CDNS_7246542145918 $T=43570 104220 0 0 $X=42600 $Y=103560
X273 2 VIA2_C_CDNS_7246542145918 $T=43570 131040 0 0 $X=42600 $Y=130380
X274 19 VIA2_C_CDNS_7246542145918 $T=107055 58225 0 0 $X=106085 $Y=57565
X275 19 VIA2_C_CDNS_7246542145918 $T=107055 85685 0 0 $X=106085 $Y=85025
X276 1 VIA2_C_CDNS_7246542145918 $T=108020 14010 0 0 $X=107050 $Y=13350
X277 1 VIA2_C_CDNS_7246542145918 $T=108020 38730 0 0 $X=107050 $Y=38070
X278 14 VIA2_C_CDNS_7246542145918 $T=109335 54665 0 0 $X=108365 $Y=54005
X279 14 VIA2_C_CDNS_7246542145918 $T=109335 87465 0 0 $X=108365 $Y=86805
X280 14 VIA2_C_CDNS_7246542145918 $T=110300 10450 0 0 $X=109330 $Y=9790
X281 14 VIA2_C_CDNS_7246542145918 $T=110300 40510 0 0 $X=109330 $Y=39850
X282 8 VIA2_C_CDNS_7246542145919 $T=5840 100660 0 0 $X=5130 $Y=100000
X283 8 VIA2_C_CDNS_7246542145919 $T=5840 134600 0 0 $X=5130 $Y=133940
X284 7 VIA2_C_CDNS_7246542145919 $T=7240 13685 0 0 $X=6530 $Y=13025
X285 7 VIA2_C_CDNS_7246542145919 $T=7240 43665 0 0 $X=6530 $Y=43005
X286 16 VIA2_C_CDNS_7246542145919 $T=9020 11905 0 0 $X=8310 $Y=11245
X287 16 VIA2_C_CDNS_7246542145919 $T=9020 41885 0 0 $X=8310 $Y=41225
X288 18 VIA2_C_CDNS_7246542145919 $T=31680 45445 0 0 $X=30970 $Y=44785
X289 17 VIA2_C_CDNS_7246542145919 $T=33460 10125 0 0 $X=32750 $Y=9465
X290 5 VIA2_C_CDNS_7246542145919 $T=45600 102440 0 0 $X=44890 $Y=101780
X291 5 VIA2_C_CDNS_7246542145919 $T=45600 136380 0 0 $X=44890 $Y=135720
X292 4 VIA2_C_CDNS_7246542145919 $T=47380 98880 0 0 $X=46670 $Y=98220
X293 4 VIA2_C_CDNS_7246542145919 $T=47380 132820 0 0 $X=46670 $Y=132160
X294 1 VIA1_C_CDNS_7246542145920 $T=95520 101635 0 0 $X=95120 $Y=100665
X295 4 VIA1_C_CDNS_7246542145920 $T=97060 99355 0 0 $X=96660 $Y=98385
X296 1 VIA1_C_CDNS_7246542145920 $T=98600 101635 0 0 $X=98200 $Y=100665
X297 4 VIA1_C_CDNS_7246542145920 $T=100140 99355 0 0 $X=99740 $Y=98385
X298 1 VIA1_C_CDNS_7246542145920 $T=101680 101635 0 0 $X=101280 $Y=100665
X299 8 VIA2_C_CDNS_7246542145927 $T=9255 74485 0 0 $X=8505 $Y=73735
X300 16 VIA2_C_CDNS_7246542145927 $T=22885 54255 0 0 $X=22135 $Y=53505
X301 10 VIA2_C_CDNS_7246542145928 $T=70110 136100 0 0 $X=68060 $Y=135350
X302 4 VIA2_C_CDNS_7246542145936 $T=118800 136695 0 0 $X=118310 $Y=134645
X303 10 VIA2_C_CDNS_7246542145936 $T=208725 98250 0 0 $X=208235 $Y=96200
X304 4 VIA1_C_CDNS_7246542145937 $T=118805 88080 0 0 $X=118315 $Y=86030
X305 4 VIA1_C_CDNS_7246542145937 $T=118805 136570 0 0 $X=118315 $Y=134520
X306 9 VIA1_C_CDNS_7246542145937 $T=208665 49725 0 0 $X=208175 $Y=47675
X307 10 VIA1_C_CDNS_7246542145937 $T=208725 98250 0 0 $X=208235 $Y=96200
X308 1 1 1 ne3_CDNS_724654214591 $T=44780 15300 0 0 $X=43980 $Y=14900
X309 1 1 1 ne3_CDNS_724654214591 $T=44780 37440 1 0 $X=43980 $Y=26870
X310 1 11 11 ne3_CDNS_724654214591 $T=51020 15300 0 0 $X=50220 $Y=14900
X311 1 11 14 ne3_CDNS_724654214591 $T=51020 37440 1 0 $X=50220 $Y=26870
X312 1 11 14 ne3_CDNS_724654214591 $T=57260 15300 0 0 $X=56460 $Y=14900
X313 1 11 11 ne3_CDNS_724654214591 $T=57260 37440 1 0 $X=56460 $Y=26870
X314 1 11 11 ne3_CDNS_724654214591 $T=63500 15300 0 0 $X=62700 $Y=14900
X315 1 11 14 ne3_CDNS_724654214591 $T=63500 37440 1 0 $X=62700 $Y=26870
X316 1 11 14 ne3_CDNS_724654214591 $T=69740 15300 0 0 $X=68940 $Y=14900
X317 1 11 11 ne3_CDNS_724654214591 $T=69740 37440 1 0 $X=68940 $Y=26870
X318 1 11 11 ne3_CDNS_724654214591 $T=75980 15300 0 0 $X=75180 $Y=14900
X319 1 11 14 ne3_CDNS_724654214591 $T=75980 37440 1 0 $X=75180 $Y=26870
X320 1 11 14 ne3_CDNS_724654214591 $T=82220 15300 0 0 $X=81420 $Y=14900
X321 1 11 11 ne3_CDNS_724654214591 $T=82220 37440 1 0 $X=81420 $Y=26870
X322 1 11 11 ne3_CDNS_724654214591 $T=88460 15300 0 0 $X=87660 $Y=14900
X323 1 11 14 ne3_CDNS_724654214591 $T=88460 37440 1 0 $X=87660 $Y=26870
X324 1 11 14 ne3_CDNS_724654214591 $T=94700 15300 0 0 $X=93900 $Y=14900
X325 1 11 11 ne3_CDNS_724654214591 $T=94700 37440 1 0 $X=93900 $Y=26870
X326 1 1 1 ne3_CDNS_724654214591 $T=100940 15300 0 0 $X=100140 $Y=14900
X327 1 1 1 ne3_CDNS_724654214591 $T=100940 37440 1 0 $X=100140 $Y=26870
X328 2 VIA1_C_CDNS_7246542145944 $T=59385 131570 0 0 $X=59245 $Y=130600
X329 12 VIA1_C_CDNS_7246542145944 $T=64925 133850 0 0 $X=64785 $Y=132880
X330 2 VIA1_C_CDNS_7246542145944 $T=65625 131570 0 0 $X=65485 $Y=130600
X331 10 VIA1_C_CDNS_7246542145944 $T=71165 136130 0 0 $X=71025 $Y=135160
X332 17 VIA1_C_CDNS_7246542145944 $T=97690 123640 0 0 $X=97550 $Y=122670
X333 13 VIA1_C_CDNS_7246542145944 $T=99230 121360 0 0 $X=99090 $Y=120390
X334 17 VIA1_C_CDNS_7246542145944 $T=99930 123640 0 0 $X=99790 $Y=122670
X335 20 VIA1_C_CDNS_7246542145944 $T=101470 119080 0 0 $X=101330 $Y=118110
X336 1 VIA2_C_CDNS_7246542145946 $T=20350 6575 0 0 $X=16220 $Y=5565
X337 1 VIA2_C_CDNS_7246542145946 $T=75360 6055 0 0 $X=71230 $Y=5045
X338 1 VIA1_C_CDNS_7246542145947 $T=20350 6575 0 0 $X=16220 $Y=5565
X339 1 VIA1_C_CDNS_7246542145947 $T=75360 6055 0 0 $X=71230 $Y=5045
X340 2 VIA1_C_CDNS_7246542145949 $T=6000 138620 0 0 $X=4210 $Y=137870
X341 2 VIA1_C_CDNS_7246542145949 $T=47220 138620 0 0 $X=45430 $Y=137870
X342 2 VIA1_C_CDNS_7246542145949 $T=59055 138620 0 0 $X=57265 $Y=137870
X343 2 VIA1_C_CDNS_7246542145949 $T=84905 138620 0 0 $X=83115 $Y=137870
X344 2 VIA1_C_CDNS_7246542145951 $T=110725 50485 0 0 $X=110235 $Y=47655
X345 2 VIA1_C_CDNS_7246542145951 $T=119195 38515 0 0 $X=118705 $Y=35685
X346 21 VIA1_C_CDNS_7246542145957 $T=296735 11275 0 0 $X=296245 $Y=7145
X347 9 VIA1_C_CDNS_7246542145957 $T=296735 36110 0 0 $X=296245 $Y=31980
X348 17 VIA2_C_CDNS_7246542145958 $T=80230 95900 0 0 $X=79480 $Y=95240
X349 21 VIA1_C_CDNS_7246542145959 $T=307595 14520 0 0 $X=307405 $Y=10480
X350 21 VIA1_C_CDNS_7246542145959 $T=307595 31270 0 0 $X=307405 $Y=27230
X351 21 VIA1_C_CDNS_7246542145959 $T=307595 48020 0 0 $X=307405 $Y=43980
X352 21 VIA1_C_CDNS_7246542145959 $T=307595 64770 0 0 $X=307405 $Y=60730
X353 21 VIA1_C_CDNS_7246542145959 $T=307595 81520 0 0 $X=307405 $Y=77480
X354 21 VIA1_C_CDNS_7246542145959 $T=307595 98270 0 0 $X=307405 $Y=94230
X355 21 VIA1_C_CDNS_7246542145959 $T=307595 115020 0 0 $X=307405 $Y=110980
X356 21 VIA1_C_CDNS_7246542145959 $T=307595 131770 0 0 $X=307405 $Y=127730
X357 21 VIA1_C_CDNS_7246542145959 $T=324350 14520 0 0 $X=324160 $Y=10480
X358 21 VIA1_C_CDNS_7246542145959 $T=324350 31270 0 0 $X=324160 $Y=27230
X359 21 VIA1_C_CDNS_7246542145959 $T=324350 48020 0 0 $X=324160 $Y=43980
X360 21 VIA1_C_CDNS_7246542145959 $T=324350 81520 0 0 $X=324160 $Y=77480
X361 21 VIA1_C_CDNS_7246542145959 $T=324350 98270 0 0 $X=324160 $Y=94230
X362 21 VIA1_C_CDNS_7246542145959 $T=324350 115020 0 0 $X=324160 $Y=110980
X363 21 VIA1_C_CDNS_7246542145959 $T=324350 131770 0 0 $X=324160 $Y=127730
X364 21 VIA1_C_CDNS_7246542145959 $T=341105 14520 0 0 $X=340915 $Y=10480
X365 21 VIA1_C_CDNS_7246542145959 $T=341105 31270 0 0 $X=340915 $Y=27230
X366 21 VIA1_C_CDNS_7246542145959 $T=341105 48020 0 0 $X=340915 $Y=43980
X367 21 VIA1_C_CDNS_7246542145959 $T=341105 64770 0 0 $X=340915 $Y=60730
X368 21 VIA1_C_CDNS_7246542145959 $T=341105 81520 0 0 $X=340915 $Y=77480
X369 21 VIA1_C_CDNS_7246542145959 $T=341105 98270 0 0 $X=340915 $Y=94230
X370 21 VIA1_C_CDNS_7246542145959 $T=341105 115020 0 0 $X=340915 $Y=110980
X371 21 VIA1_C_CDNS_7246542145959 $T=341105 131770 0 0 $X=340915 $Y=127730
X372 21 VIA1_C_CDNS_7246542145959 $T=357860 14520 0 0 $X=357670 $Y=10480
X373 21 VIA1_C_CDNS_7246542145959 $T=357860 31270 0 0 $X=357670 $Y=27230
X374 21 VIA1_C_CDNS_7246542145959 $T=357860 48020 0 0 $X=357670 $Y=43980
X375 21 VIA1_C_CDNS_7246542145959 $T=357860 64770 0 0 $X=357670 $Y=60730
X376 21 VIA1_C_CDNS_7246542145959 $T=357860 81520 0 0 $X=357670 $Y=77480
X377 21 VIA1_C_CDNS_7246542145959 $T=357860 98270 0 0 $X=357670 $Y=94230
X378 21 VIA1_C_CDNS_7246542145959 $T=357860 115020 0 0 $X=357670 $Y=110980
X379 21 VIA1_C_CDNS_7246542145959 $T=357860 131770 0 0 $X=357670 $Y=127730
X380 8 6 6 2 1 pe3_CDNS_7246542145911 $T=9635 78185 0 0 $X=8125 $Y=77155
X381 5 6 19 2 1 pe3_CDNS_7246542145911 $T=23440 78185 0 0 $X=21930 $Y=77155
X382 7 3 3 1 ne3_CDNS_7246542145912 $T=10345 55405 0 0 $X=9545 $Y=55005
X383 16 3 6 1 ne3_CDNS_7246542145912 $T=22730 55545 0 0 $X=21930 $Y=55145
X384 1 14 4 1 ne3_CDNS_7246542145912 $T=95790 103175 0 0 $X=94990 $Y=102775
X385 9 21 1 rpp1k1_3_CDNS_7246542145913 $T=287735 7255 1 180 $X=159445 $Y=7035
X386 4 22 1 rpp1k1_3_CDNS_7246542145914 $T=123895 47740 0 0 $X=118735 $Y=47520
X387 1 1 1 1 ne3_CDNS_7246542145915 $T=13130 16755 0 0 $X=12330 $Y=16355
X388 1 1 1 1 ne3_CDNS_7246542145915 $T=13130 38815 1 0 $X=12330 $Y=28245
X389 1 7 16 1 ne3_CDNS_7246542145915 $T=15370 16755 0 0 $X=14570 $Y=16355
X390 1 7 7 1 ne3_CDNS_7246542145915 $T=15370 38815 1 0 $X=14570 $Y=28245
X391 1 7 7 1 ne3_CDNS_7246542145915 $T=17610 16755 0 0 $X=16810 $Y=16355
X392 1 7 16 1 ne3_CDNS_7246542145915 $T=17610 38815 1 0 $X=16810 $Y=28245
X393 1 7 17 1 ne3_CDNS_7246542145915 $T=19850 16755 0 0 $X=19050 $Y=16355
X394 1 7 18 1 ne3_CDNS_7246542145915 $T=19850 38815 1 0 $X=19050 $Y=28245
X395 1 7 16 1 ne3_CDNS_7246542145915 $T=22090 16755 0 0 $X=21290 $Y=16355
X396 1 7 7 1 ne3_CDNS_7246542145915 $T=22090 38815 1 0 $X=21290 $Y=28245
X397 1 7 7 1 ne3_CDNS_7246542145915 $T=24330 16755 0 0 $X=23530 $Y=16355
X398 1 7 16 1 ne3_CDNS_7246542145915 $T=24330 38815 1 0 $X=23530 $Y=28245
X399 1 1 1 1 ne3_CDNS_7246542145915 $T=26570 16755 0 0 $X=25770 $Y=16355
X400 1 1 1 1 ne3_CDNS_7246542145915 $T=26570 38815 1 0 $X=25770 $Y=28245
X401 17 4 13 1 ne3_CDNS_7246542145915 $T=97960 125180 0 0 $X=97160 $Y=124780
X402 17 15 20 1 ne3_CDNS_7246542145915 $T=100200 125180 0 0 $X=99400 $Y=124780
X403 19 19 19 2 1 pe3_CDNS_7246542145916 $T=43105 60145 0 0 $X=41595 $Y=59115
X404 19 19 19 2 1 pe3_CDNS_7246542145916 $T=43105 83765 1 0 $X=41595 $Y=72735
X405 19 10 14 2 1 pe3_CDNS_7246542145916 $T=49345 60145 0 0 $X=47835 $Y=59115
X406 19 9 11 2 1 pe3_CDNS_7246542145916 $T=49345 83765 1 0 $X=47835 $Y=72735
X407 19 9 11 2 1 pe3_CDNS_7246542145916 $T=55585 60145 0 0 $X=54075 $Y=59115
X408 19 10 14 2 1 pe3_CDNS_7246542145916 $T=55585 83765 1 0 $X=54075 $Y=72735
X409 2 12 12 2 1 pe3_CDNS_7246542145916 $T=59655 129400 1 0 $X=58145 $Y=118370
X410 19 10 14 2 1 pe3_CDNS_7246542145916 $T=61825 60145 0 0 $X=60315 $Y=59115
X411 19 9 11 2 1 pe3_CDNS_7246542145916 $T=61825 83765 1 0 $X=60315 $Y=72735
X412 2 12 10 2 1 pe3_CDNS_7246542145916 $T=65895 129400 1 0 $X=64385 $Y=118370
X413 19 9 11 2 1 pe3_CDNS_7246542145916 $T=68065 60145 0 0 $X=66555 $Y=59115
X414 19 10 14 2 1 pe3_CDNS_7246542145916 $T=68065 83765 1 0 $X=66555 $Y=72735
X415 19 10 14 2 1 pe3_CDNS_7246542145916 $T=74305 60145 0 0 $X=72795 $Y=59115
X416 19 9 11 2 1 pe3_CDNS_7246542145916 $T=74305 83765 1 0 $X=72795 $Y=72735
X417 2 13 13 2 1 pe3_CDNS_7246542145916 $T=79075 125320 0 0 $X=77565 $Y=124290
X418 19 9 11 2 1 pe3_CDNS_7246542145916 $T=80545 60145 0 0 $X=79035 $Y=59115
X419 19 10 14 2 1 pe3_CDNS_7246542145916 $T=80545 83765 1 0 $X=79035 $Y=72735
X420 2 13 20 2 1 pe3_CDNS_7246542145916 $T=85315 125320 0 0 $X=83805 $Y=124290
X421 19 10 14 2 1 pe3_CDNS_7246542145916 $T=86785 60145 0 0 $X=85275 $Y=59115
X422 19 9 11 2 1 pe3_CDNS_7246542145916 $T=86785 83765 1 0 $X=85275 $Y=72735
X423 19 9 11 2 1 pe3_CDNS_7246542145916 $T=93025 60145 0 0 $X=91515 $Y=59115
X424 19 10 14 2 1 pe3_CDNS_7246542145916 $T=93025 83765 1 0 $X=91515 $Y=72735
X425 19 19 19 2 1 pe3_CDNS_7246542145916 $T=99265 60145 0 0 $X=97755 $Y=59115
X426 19 19 19 2 1 pe3_CDNS_7246542145916 $T=99265 83765 1 0 $X=97755 $Y=72735
X427 12 20 18 2 1 pe3_CDNS_7246542145917 $T=62750 104210 0 0 $X=61240 $Y=103180
X428 1 15 1 ne3_CDNS_7246542145918 $T=110195 126990 0 0 $X=109395 $Y=126590
X429 15 23 1 ne3_CDNS_7246542145918 $T=110195 130510 0 0 $X=109395 $Y=130110
X430 23 2 1 ne3_CDNS_7246542145918 $T=110195 134045 0 0 $X=109395 $Y=133645
X431 2 2 2 1 pe3_CDNS_7246542145919 $T=10660 106140 0 0 $X=9150 $Y=105110
X432 2 2 2 1 pe3_CDNS_7246542145919 $T=10660 129120 1 0 $X=9150 $Y=118090
X433 2 8 4 1 pe3_CDNS_7246542145919 $T=12900 106140 0 0 $X=11390 $Y=105110
X434 2 8 4 1 pe3_CDNS_7246542145919 $T=12900 129120 1 0 $X=11390 $Y=118090
X435 2 8 4 1 pe3_CDNS_7246542145919 $T=15140 106140 0 0 $X=13630 $Y=105110
X436 2 8 4 1 pe3_CDNS_7246542145919 $T=15140 129120 1 0 $X=13630 $Y=118090
X437 2 8 5 1 pe3_CDNS_7246542145919 $T=17380 106140 0 0 $X=15870 $Y=105110
X438 2 8 8 1 pe3_CDNS_7246542145919 $T=17380 129120 1 0 $X=15870 $Y=118090
X439 2 8 4 1 pe3_CDNS_7246542145919 $T=19620 106140 0 0 $X=18110 $Y=105110
X440 2 8 4 1 pe3_CDNS_7246542145919 $T=19620 129120 1 0 $X=18110 $Y=118090
X441 2 8 4 1 pe3_CDNS_7246542145919 $T=21860 106140 0 0 $X=20350 $Y=105110
X442 2 8 4 1 pe3_CDNS_7246542145919 $T=21860 129120 1 0 $X=20350 $Y=118090
X443 2 8 8 1 pe3_CDNS_7246542145919 $T=24100 106140 0 0 $X=22590 $Y=105110
X444 2 8 5 1 pe3_CDNS_7246542145919 $T=24100 129120 1 0 $X=22590 $Y=118090
X445 2 8 5 1 pe3_CDNS_7246542145919 $T=26340 106140 0 0 $X=24830 $Y=105110
X446 2 8 8 1 pe3_CDNS_7246542145919 $T=26340 129120 1 0 $X=24830 $Y=118090
X447 2 8 4 1 pe3_CDNS_7246542145919 $T=28580 106140 0 0 $X=27070 $Y=105110
X448 2 8 4 1 pe3_CDNS_7246542145919 $T=28580 129120 1 0 $X=27070 $Y=118090
X449 2 8 4 1 pe3_CDNS_7246542145919 $T=30820 106140 0 0 $X=29310 $Y=105110
X450 2 8 4 1 pe3_CDNS_7246542145919 $T=30820 129120 1 0 $X=29310 $Y=118090
X451 2 8 8 1 pe3_CDNS_7246542145919 $T=33060 106140 0 0 $X=31550 $Y=105110
X452 2 8 5 1 pe3_CDNS_7246542145919 $T=33060 129120 1 0 $X=31550 $Y=118090
X453 2 8 4 1 pe3_CDNS_7246542145919 $T=35300 106140 0 0 $X=33790 $Y=105110
X454 2 8 4 1 pe3_CDNS_7246542145919 $T=35300 129120 1 0 $X=33790 $Y=118090
X455 2 8 4 1 pe3_CDNS_7246542145919 $T=37540 106140 0 0 $X=36030 $Y=105110
X456 2 8 4 1 pe3_CDNS_7246542145919 $T=37540 129120 1 0 $X=36030 $Y=118090
X457 2 2 2 1 pe3_CDNS_7246542145919 $T=39780 106140 0 0 $X=38270 $Y=105110
X458 2 2 2 1 pe3_CDNS_7246542145919 $T=39780 129120 1 0 $X=38270 $Y=118090
X459 4 24 1 rpp1k1_3_CDNS_7246542145920 $T=123895 96235 0 0 $X=118735 $Y=96015
X460 22 9 1 rpp1k1_3_CDNS_7246542145920 $T=213685 47740 0 0 $X=208525 $Y=47520
X461 24 10 1 rpp1k1_3_CDNS_7246542145920 $T=213685 96235 0 0 $X=208525 $Y=96015
Q0 1 1 21 qpvc3 $X=302595 $Y=9520 $dt=4
Q1 1 1 21 qpvc3 $X=302595 $Y=26270 $dt=4
Q2 1 1 21 qpvc3 $X=302595 $Y=43020 $dt=4
Q3 1 1 21 qpvc3 $X=302595 $Y=59770 $dt=4
Q4 1 1 21 qpvc3 $X=302595 $Y=76520 $dt=4
Q5 1 1 21 qpvc3 $X=302595 $Y=93270 $dt=4
Q6 1 1 21 qpvc3 $X=302595 $Y=110020 $dt=4
Q7 1 1 21 qpvc3 $X=302595 $Y=126770 $dt=4
Q8 1 1 21 qpvc3 $X=319350 $Y=9520 $dt=4
Q9 1 1 21 qpvc3 $X=319350 $Y=26270 $dt=4
Q10 1 1 21 qpvc3 $X=319350 $Y=43020 $dt=4
Q11 1 1 10 qpvc3 $X=319350 $Y=59770 $dt=4
Q12 1 1 21 qpvc3 $X=319350 $Y=76520 $dt=4
Q13 1 1 21 qpvc3 $X=319350 $Y=93270 $dt=4
Q14 1 1 21 qpvc3 $X=319350 $Y=110020 $dt=4
Q15 1 1 21 qpvc3 $X=319350 $Y=126770 $dt=4
Q16 1 1 21 qpvc3 $X=336105 $Y=9520 $dt=4
Q17 1 1 21 qpvc3 $X=336105 $Y=26270 $dt=4
Q18 1 1 21 qpvc3 $X=336105 $Y=43020 $dt=4
Q19 1 1 21 qpvc3 $X=336105 $Y=59770 $dt=4
Q20 1 1 21 qpvc3 $X=336105 $Y=76520 $dt=4
Q21 1 1 21 qpvc3 $X=336105 $Y=93270 $dt=4
Q22 1 1 21 qpvc3 $X=336105 $Y=110020 $dt=4
Q23 1 1 21 qpvc3 $X=336105 $Y=126770 $dt=4
Q24 1 1 21 qpvc3 $X=352860 $Y=9520 $dt=4
Q25 1 1 21 qpvc3 $X=352860 $Y=26270 $dt=4
Q26 1 1 21 qpvc3 $X=352860 $Y=43020 $dt=4
Q27 1 1 21 qpvc3 $X=352860 $Y=59770 $dt=4
Q28 1 1 21 qpvc3 $X=352860 $Y=76520 $dt=4
Q29 1 1 21 qpvc3 $X=352860 $Y=93270 $dt=4
Q30 1 1 21 qpvc3 $X=352860 $Y=110020 $dt=4
Q31 1 1 21 qpvc3 $X=352860 $Y=126770 $dt=4
D32 1 2 p_dnw AREA=1.07147e-09 PJ=0.0001732 perimeter=0.0001732 $X=3950 $Y=96990 $dt=5
D33 1 2 p_dnw AREA=2.50005e-10 PJ=8.653e-05 perimeter=8.653e-05 $X=6985 $Y=72595 $dt=5
D34 1 2 p_dnw AREA=1.35123e-09 PJ=0.00022788 perimeter=0.00022788 $X=35895 $Y=52775 $dt=5
D35 1 2 p_dnw AREA=3.30547e-10 PJ=0.00010554 perimeter=0.00010554 $X=57005 $Y=102040 $dt=5
D36 1 2 p_dnw AREA=1.64117e-10 PJ=7.372e-05 perimeter=7.372e-05 $X=76425 $Y=117950 $dt=5
D37 1 2 p_dnw AREA=1.17512e-09 PJ=0.00013712 perimeter=0.00013712 $X=119255 $Y=7325 $dt=5
D38 1 2 p_dnw3 AREA=3.99668e-10 PJ=0 perimeter=0 $X=9150 $Y=105110 $dt=8
D39 1 2 p_dnw3 AREA=3.99668e-10 PJ=0 perimeter=0 $X=9150 $Y=118090 $dt=8
D40 1 2 p_dnw3 AREA=7.74011e-10 PJ=0 perimeter=0 $X=41595 $Y=59115 $dt=8
D41 1 2 p_dnw3 AREA=7.74011e-10 PJ=0 perimeter=0 $X=41595 $Y=72735 $dt=8
D42 1 2 p_dnw3 AREA=1.71976e-10 PJ=0 perimeter=0 $X=58145 $Y=118370 $dt=8
D43 1 2 p_dnw3 AREA=1.71976e-10 PJ=0 perimeter=0 $X=77565 $Y=124290 $dt=8
C44 14 4 area=9e-10 perimeter=0.00012 $[cmm5t] $X=121395 $Y=9465 $dt=11
.ends bandgap_su

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: mosvc3_CDNS_7246542145921                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt mosvc3_CDNS_7246542145921 1 2
** N=2 EP=2 FDC=2
X0 2 1 1 MOSVC3 w=2.5e-05 l=3e-05 $X=0 $Y=0 $dt=3
D1 1 1 p_dnw3 AREA=6.7176e-11 PJ=0.00011492 perimeter=0.00011492 $X=-800 $Y=-430 $dt=8
.ends mosvc3_CDNS_7246542145921

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246542145966                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246542145966 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246542145966

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246542145968                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246542145968 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246542145968

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246542145972                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246542145972 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246542145972

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246542145973                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246542145973 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246542145973

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246542145977                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246542145977 1 2
** N=2 EP=2 FDC=0
.ends VIA2_C_CDNS_7246542145977

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3i_6_CDNS_7246542145922                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3i_6_CDNS_7246542145922 1 2 3
** N=3 EP=3 FDC=4
X0 1 3 3 1 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=4.8e-12 ps=1.054e-05 pd=2.096e-05 $X=0 $Y=0 $dt=2
X1 3 3 1 1 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=4.8e-12 ad=2.7e-12 ps=2.096e-05 pd=1.054e-05 $X=3040 $Y=0 $dt=2
D2 1 2 p_ddnw AREA=3.07331e-10 PJ=7.576e-05 perimeter=7.576e-05 $X=-6110 $Y=-4940 $dt=6
D3 1 2 p_dipdnwmv AREA=7.49452e-11 PJ=4.496e-05 perimeter=4.496e-05 $X=-2260 $Y=-1090 $dt=7
.ends ne3i_6_CDNS_7246542145922

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246542145923                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246542145923 1 2 3
** N=3 EP=3 FDC=2
M0 2 2 1 1 pe3 L=1e-05 W=2e-06 AD=9.6e-13 AS=9.6e-13 PD=4.96e-06 PS=4.96e-06 $X=0 $Y=0 $dt=1
D1 3 1 p_dnw3 AREA=4.57434e-11 PJ=3.138e-05 perimeter=3.138e-05 $X=-910 $Y=-1440 $dt=8
.ends pe3_CDNS_7246542145923

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7246542145924                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7246542145924 1 2 3 4
** N=4 EP=4 FDC=2
M0 3 2 1 4 ne3 L=2.5e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
M1 1 2 3 4 ne3 L=2.5e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=3040 $Y=0 $dt=0
.ends ne3_CDNS_7246542145924

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246542145925                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246542145925 1 2 3 4 5
** N=5 EP=5 FDC=3
M0 3 2 1 4 pe3 L=2.5e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=2.5e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=3040 $Y=0 $dt=1
D2 5 4 p_dnw3 AREA=1.03234e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=8
.ends pe3_CDNS_7246542145925

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246542145926                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246542145926 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 3 2 1 4 pe3 L=2.5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
D1 5 4 p_dnw3 AREA=6.65712e-11 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=8
.ends pe3_CDNS_7246542145926

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246542145927                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246542145927 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
M0 3 2 1 1 pe3 L=2.5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_7246542145927

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3i_6_CDNS_7246542145928                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3i_6_CDNS_7246542145928 1 2 3 4 5
** N=5 EP=5 FDC=10
X0 3 4 5 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=4.8e-12 ps=1.054e-05 pd=2.096e-05 $X=0 $Y=0 $dt=2
X1 5 4 3 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=2.7e-12 ps=1.054e-05 pd=1.054e-05 $X=3040 $Y=0 $dt=2
X2 3 4 5 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=2.7e-12 ps=1.054e-05 pd=1.054e-05 $X=6080 $Y=0 $dt=2
X3 5 4 3 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=2.7e-12 ps=1.054e-05 pd=1.054e-05 $X=9120 $Y=0 $dt=2
X4 3 4 5 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=2.7e-12 ps=1.054e-05 pd=1.054e-05 $X=12160 $Y=0 $dt=2
X5 5 4 3 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=2.7e-12 ps=1.054e-05 pd=1.054e-05 $X=15200 $Y=0 $dt=2
X6 3 4 5 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=2.7e-12 ps=1.054e-05 pd=1.054e-05 $X=18240 $Y=0 $dt=2
X7 5 4 3 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=4.8e-12 ad=2.7e-12 ps=2.096e-05 pd=1.054e-05 $X=21280 $Y=0 $dt=2
D8 1 2 p_ddnw AREA=5.2432e-10 PJ=0.00011224 perimeter=0.00011224 $X=-6110 $Y=-4940 $dt=6
D9 3 2 p_dipdnwmv AREA=1.51486e-10 PJ=8.144e-05 perimeter=8.144e-05 $X=-2260 $Y=-1090 $dt=7
.ends ne3i_6_CDNS_7246542145928

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7246542145929                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7246542145929 1 2 3
*.DEVICECLIMB
** N=3 EP=3 FDC=1
R0 2 1 L=0.0002878 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=10
.ends rpp1k1_3_CDNS_7246542145929

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: constant_gm                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt constant_gm 1 2 3 4 5
** N=16 EP=5 FDC=56
X0 6 VIA2_C_CDNS_724654214593 $T=14445 92470 0 0 $X=13735 $Y=92070
X1 6 VIA2_C_CDNS_724654214593 $T=14445 111830 0 0 $X=13735 $Y=111430
X2 7 VIA2_C_CDNS_724654214593 $T=48025 75790 0 0 $X=47315 $Y=75390
X3 7 VIA2_C_CDNS_724654214593 $T=48025 91190 0 0 $X=47315 $Y=90790
X4 7 VIA2_C_CDNS_724654214593 $T=48025 110550 0 0 $X=47315 $Y=110150
X5 8 VIA2_C_CDNS_724654214593 $T=49805 93750 0 0 $X=49095 $Y=93350
X6 8 VIA2_C_CDNS_724654214593 $T=49805 113110 0 0 $X=49095 $Y=112710
X7 9 VIA2_C_CDNS_724654214593 $T=51585 95030 0 0 $X=50875 $Y=94630
X8 9 VIA2_C_CDNS_724654214593 $T=51585 114390 0 0 $X=50875 $Y=113990
X9 10 VIA2_C_CDNS_724654214593 $T=53365 115670 0 0 $X=52655 $Y=115270
X10 7 VIA1_C_CDNS_724654214594 $T=23755 75790 0 0 $X=23615 $Y=75340
X11 7 VIA1_C_CDNS_724654214594 $T=23755 91190 0 0 $X=23615 $Y=90740
X12 7 VIA1_C_CDNS_724654214594 $T=27495 75790 0 0 $X=27355 $Y=75340
X13 7 VIA1_C_CDNS_724654214594 $T=27495 91190 0 0 $X=27355 $Y=90740
X14 7 VIA1_C_CDNS_724654214594 $T=31235 75790 0 0 $X=31095 $Y=75340
X15 7 VIA1_C_CDNS_724654214594 $T=31235 91190 0 0 $X=31095 $Y=90740
X16 7 VIA1_C_CDNS_724654214594 $T=34975 75790 0 0 $X=34835 $Y=75340
X17 7 VIA1_C_CDNS_724654214594 $T=34975 91190 0 0 $X=34835 $Y=90740
X18 7 VIA1_C_CDNS_724654214594 $T=38715 91190 0 0 $X=38575 $Y=90740
X19 11 VIA1_C_CDNS_7246542145911 $T=12910 70305 0 0 $X=11990 $Y=70115
X20 11 VIA1_C_CDNS_7246542145911 $T=15950 70305 0 0 $X=15030 $Y=70115
X21 11 VIA1_C_CDNS_7246542145911 $T=23060 70305 0 0 $X=22140 $Y=70115
X22 11 VIA1_C_CDNS_7246542145911 $T=26100 70305 0 0 $X=25180 $Y=70115
X23 12 VIA1_C_CDNS_7246542145911 $T=26710 50605 0 0 $X=25790 $Y=50415
X24 12 VIA1_C_CDNS_7246542145911 $T=29750 50605 0 0 $X=28830 $Y=50415
X25 11 VIA1_C_CDNS_7246542145911 $T=33815 70305 0 0 $X=32895 $Y=70115
X26 12 VIA1_C_CDNS_7246542145911 $T=36040 50605 0 0 $X=35120 $Y=50415
X27 11 VIA1_C_CDNS_7246542145911 $T=36855 70305 0 0 $X=35935 $Y=70115
X28 12 VIA1_C_CDNS_7246542145911 $T=39080 50605 0 0 $X=38160 $Y=50415
X29 11 VIA1_C_CDNS_7246542145911 $T=44630 70305 0 0 $X=43710 $Y=70115
X30 11 VIA1_C_CDNS_7246542145911 $T=47670 70305 0 0 $X=46750 $Y=70115
X31 2 VIA1_C_CDNS_7246542145912 $T=18495 89660 0 0 $X=18355 $Y=88950
X32 2 VIA1_C_CDNS_7246542145912 $T=18495 109020 0 0 $X=18355 $Y=108310
X33 2 VIA1_C_CDNS_7246542145912 $T=21535 89660 0 0 $X=21395 $Y=88950
X34 2 VIA1_C_CDNS_7246542145912 $T=21535 109020 0 0 $X=21395 $Y=108310
X35 2 VIA1_C_CDNS_7246542145912 $T=22235 89660 0 0 $X=22095 $Y=88950
X36 2 VIA1_C_CDNS_7246542145912 $T=22235 109020 0 0 $X=22095 $Y=108310
X37 2 VIA1_C_CDNS_7246542145912 $T=25975 89660 0 0 $X=25835 $Y=88950
X38 2 VIA1_C_CDNS_7246542145912 $T=25975 109020 0 0 $X=25835 $Y=108310
X39 2 VIA1_C_CDNS_7246542145912 $T=29715 89660 0 0 $X=29575 $Y=88950
X40 2 VIA1_C_CDNS_7246542145912 $T=29715 109020 0 0 $X=29575 $Y=108310
X41 2 VIA1_C_CDNS_7246542145912 $T=33455 89660 0 0 $X=33315 $Y=88950
X42 2 VIA1_C_CDNS_7246542145912 $T=33455 109020 0 0 $X=33315 $Y=108310
X43 2 VIA1_C_CDNS_7246542145912 $T=37195 89660 0 0 $X=37055 $Y=88950
X44 2 VIA1_C_CDNS_7246542145912 $T=37195 109020 0 0 $X=37055 $Y=108310
X45 2 VIA1_C_CDNS_7246542145912 $T=40235 89660 0 0 $X=40095 $Y=88950
X46 2 VIA1_C_CDNS_7246542145912 $T=40935 89660 0 0 $X=40795 $Y=88950
X47 2 VIA1_C_CDNS_7246542145912 $T=40935 109020 0 0 $X=40795 $Y=108310
X48 2 VIA1_C_CDNS_7246542145912 $T=43975 89660 0 0 $X=43835 $Y=88950
X49 2 VIA1_C_CDNS_7246542145912 $T=43975 109020 0 0 $X=43835 $Y=108310
X50 2 VIA2_C_CDNS_7246542145919 $T=16225 89660 0 0 $X=15515 $Y=89000
X51 2 VIA2_C_CDNS_7246542145919 $T=16225 109020 0 0 $X=15515 $Y=108360
X52 2 VIA2_C_CDNS_7246542145919 $T=46245 89660 0 0 $X=45535 $Y=89000
X53 2 VIA2_C_CDNS_7246542145919 $T=46245 109020 0 0 $X=45535 $Y=108360
X54 9 VIA2_C_CDNS_7246542145927 $T=51305 66015 0 0 $X=50555 $Y=65265
X55 1 VIA1_C_CDNS_7246542145949 $T=20695 3535 0 0 $X=18905 $Y=2785
X56 6 VIA2_C_CDNS_7246542145958 $T=19200 68420 0 0 $X=18450 $Y=67760
X57 7 VIA2_C_CDNS_7246542145958 $T=29865 68705 0 0 $X=29115 $Y=68045
X58 8 VIA2_C_CDNS_7246542145958 $T=40615 68490 0 0 $X=39865 $Y=67830
X59 6 VIA1_C_CDNS_7246542145966 $T=11390 57075 0 0 $X=10990 $Y=56625
X60 12 VIA1_C_CDNS_7246542145966 $T=14430 55795 0 0 $X=14030 $Y=55345
X61 6 VIA1_C_CDNS_7246542145966 $T=17470 57075 0 0 $X=17070 $Y=56625
X62 7 VIA1_C_CDNS_7246542145966 $T=21540 55655 0 0 $X=21140 $Y=55205
X63 11 VIA1_C_CDNS_7246542145966 $T=24580 56935 0 0 $X=24180 $Y=56485
X64 13 VIA1_C_CDNS_7246542145966 $T=25190 37045 0 0 $X=24790 $Y=36595
X65 9 VIA1_C_CDNS_7246542145966 $T=25275 95030 0 0 $X=24875 $Y=94580
X66 9 VIA1_C_CDNS_7246542145966 $T=25275 114390 0 0 $X=24875 $Y=113940
X67 7 VIA1_C_CDNS_7246542145966 $T=27620 55655 0 0 $X=27220 $Y=55205
X68 12 VIA1_C_CDNS_7246542145966 $T=28230 38325 0 0 $X=27830 $Y=37875
X69 6 VIA1_C_CDNS_7246542145966 $T=29015 111830 0 0 $X=28615 $Y=111380
X70 13 VIA1_C_CDNS_7246542145966 $T=31270 37045 0 0 $X=30870 $Y=36595
X71 8 VIA1_C_CDNS_7246542145966 $T=32295 55655 0 0 $X=31895 $Y=55205
X72 6 VIA1_C_CDNS_7246542145966 $T=32755 92470 0 0 $X=32355 $Y=92020
X73 14 VIA1_C_CDNS_7246542145966 $T=34520 37045 0 0 $X=34120 $Y=36595
X74 3 VIA1_C_CDNS_7246542145966 $T=35335 56935 0 0 $X=34935 $Y=56485
X75 8 VIA1_C_CDNS_7246542145966 $T=36495 93750 0 0 $X=36095 $Y=93300
X76 8 VIA1_C_CDNS_7246542145966 $T=36495 113110 0 0 $X=36095 $Y=112660
X77 11 VIA1_C_CDNS_7246542145966 $T=37560 38325 0 0 $X=37160 $Y=37875
X78 8 VIA1_C_CDNS_7246542145966 $T=38375 55655 0 0 $X=37975 $Y=55205
X79 10 VIA1_C_CDNS_7246542145966 $T=40235 115670 0 0 $X=39835 $Y=115220
X80 14 VIA1_C_CDNS_7246542145966 $T=40600 37045 0 0 $X=40200 $Y=36595
X81 9 VIA1_C_CDNS_7246542145966 $T=43110 55655 0 0 $X=42710 $Y=55205
X82 4 VIA1_C_CDNS_7246542145966 $T=46150 56935 0 0 $X=45750 $Y=56485
X83 9 VIA1_C_CDNS_7246542145966 $T=49190 55655 0 0 $X=48790 $Y=55205
X84 15 VIA1_C_CDNS_7246542145968 $T=64765 41965 0 0 $X=62975 $Y=41475
X85 1 VIA1_C_CDNS_7246542145968 $T=77600 41965 0 0 $X=75810 $Y=41475
X86 1 VIA1_C_CDNS_7246542145968 $T=77650 33280 0 0 $X=75860 $Y=32790
X87 3 VIA2_C_CDNS_7246542145972 $T=35335 56935 0 0 $X=33805 $Y=56445
X88 14 VIA2_C_CDNS_7246542145972 $T=36610 37055 0 0 $X=35080 $Y=36565
X89 4 VIA2_C_CDNS_7246542145972 $T=46150 56935 0 0 $X=44620 $Y=56445
X90 7 VIA1_C_CDNS_7246542145973 $T=29015 91190 0 0 $X=28045 $Y=91050
X91 7 VIA1_C_CDNS_7246542145973 $T=32755 110550 0 0 $X=31785 $Y=110410
X92 2 1 VIA2_C_CDNS_7246542145977 $T=16225 120015 0 0 $X=14695 $Y=118485
X93 2 1 VIA2_C_CDNS_7246542145977 $T=46240 119870 0 0 $X=44710 $Y=118340
X94 1 2 13 ne3i_6_CDNS_7246542145922 $T=18020 14875 0 0 $X=7250 $Y=5275
X95 16 12 1 pe3_CDNS_7246542145923 $T=10155 41775 0 0 $X=8645 $Y=39735
X96 11 16 1 pe3_CDNS_7246542145923 $T=20155 47905 1 180 $X=8645 $Y=45865
X97 13 12 12 1 ne3_CDNS_7246542145924 $T=25460 39505 0 0 $X=24660 $Y=39105
X98 14 12 11 1 ne3_CDNS_7246542145924 $T=34790 39505 0 0 $X=33990 $Y=39105
X99 6 11 12 2 1 pe3_CDNS_7246542145925 $T=11660 58745 0 0 $X=10150 $Y=57715
X100 7 11 11 2 1 pe3_CDNS_7246542145925 $T=21810 58745 0 0 $X=20300 $Y=57715
X101 8 11 3 2 1 pe3_CDNS_7246542145925 $T=32565 58745 0 0 $X=31055 $Y=57715
X102 9 11 4 2 1 pe3_CDNS_7246542145925 $T=43380 58745 0 0 $X=41870 $Y=57715
X103 10 11 5 2 1 pe3_CDNS_7246542145926 $T=53845 58745 0 0 $X=52335 $Y=57715
X104 2 2 2 1 pe3_CDNS_7246542145927 $T=18765 87600 1 0 $X=17255 $Y=76570
X105 2 2 2 1 pe3_CDNS_7246542145927 $T=18765 106960 1 0 $X=17255 $Y=95930
X106 2 7 9 1 pe3_CDNS_7246542145927 $T=22505 87600 1 0 $X=20995 $Y=76570
X107 2 7 9 1 pe3_CDNS_7246542145927 $T=22505 106960 1 0 $X=20995 $Y=95930
X108 2 7 7 1 pe3_CDNS_7246542145927 $T=26245 87600 1 0 $X=24735 $Y=76570
X109 2 7 6 1 pe3_CDNS_7246542145927 $T=26245 106960 1 0 $X=24735 $Y=95930
X110 2 7 6 1 pe3_CDNS_7246542145927 $T=29985 87600 1 0 $X=28475 $Y=76570
X111 2 7 7 1 pe3_CDNS_7246542145927 $T=29985 106960 1 0 $X=28475 $Y=95930
X112 2 7 8 1 pe3_CDNS_7246542145927 $T=33725 87600 1 0 $X=32215 $Y=76570
X113 2 7 8 1 pe3_CDNS_7246542145927 $T=33725 106960 1 0 $X=32215 $Y=95930
X114 2 2 2 1 pe3_CDNS_7246542145927 $T=37465 87600 1 0 $X=35955 $Y=76570
X115 2 7 10 1 pe3_CDNS_7246542145927 $T=37465 106960 1 0 $X=35955 $Y=95930
X116 2 2 2 1 pe3_CDNS_7246542145927 $T=41205 87600 1 0 $X=39695 $Y=76570
X117 2 2 2 1 pe3_CDNS_7246542145927 $T=41205 106960 1 0 $X=39695 $Y=95930
X118 1 2 15 13 14 ne3i_6_CDNS_7246542145928 $T=48275 14875 0 0 $X=37505 $Y=5275
X119 1 15 2 rpp1k1_3_CDNS_7246542145929 $T=62765 46455 1 90 $X=62545 $Y=41295
D0 1 2 p_dnw AREA=4.77568e-10 PJ=0.00014131 perimeter=0.00014131 $X=7700 $Y=53605 $dt=5
D1 1 2 p_dnw AREA=1.16854e-09 PJ=0.00017172 perimeter=0.00017172 $X=12555 $Y=74150 $dt=5
D2 1 2 p_dnw AREA=1.48411e-09 PJ=0.00019385 perimeter=0.00019385 $X=61625 $Y=40375 $dt=5
D3 1 2 p_dnw3 AREA=3.37198e-10 PJ=0 perimeter=0 $X=17255 $Y=76570 $dt=8
D4 1 2 p_dnw3 AREA=3.37198e-10 PJ=0 perimeter=0 $X=17255 $Y=95930 $dt=8
.ends constant_gm

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: bias                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt bias 7 6 5 9 2 4 3
** N=9 EP=7 FDC=460
X0 1 VIA2_C_CDNS_724654214590 $T=474425 51395 0 0 $X=473675 $Y=50645
X1 2 3 1 4 5 6 7 ref_bias $T=469540 4625 0 0 $X=471000 $Y=6590
X2 2 3 8 7 bandgap_su $T=97685 3355 0 0 $X=99220 $Y=6370
X3 2 3 mosvc3_CDNS_7246542145921 $T=25775 183420 1 0 $X=24975 $Y=157800
X4 2 3 mosvc3_CDNS_7246542145921 $T=25775 185680 0 0 $X=24975 $Y=185250
X5 2 3 mosvc3_CDNS_7246542145921 $T=58775 183420 1 0 $X=57975 $Y=157800
X6 2 3 mosvc3_CDNS_7246542145921 $T=58775 185680 0 0 $X=57975 $Y=185250
X7 2 3 mosvc3_CDNS_7246542145921 $T=91775 183420 1 0 $X=90975 $Y=157800
X8 2 3 mosvc3_CDNS_7246542145921 $T=91775 185680 0 0 $X=90975 $Y=185250
X9 2 3 mosvc3_CDNS_7246542145921 $T=124775 183420 1 0 $X=123975 $Y=157800
X10 2 3 mosvc3_CDNS_7246542145921 $T=124775 185680 0 0 $X=123975 $Y=185250
X11 2 3 mosvc3_CDNS_7246542145921 $T=157775 183420 1 0 $X=156975 $Y=157800
X12 2 3 mosvc3_CDNS_7246542145921 $T=157775 185680 0 0 $X=156975 $Y=185250
X13 2 3 mosvc3_CDNS_7246542145921 $T=190775 183420 1 0 $X=189975 $Y=157800
X14 2 3 mosvc3_CDNS_7246542145921 $T=190775 185680 0 0 $X=189975 $Y=185250
X15 2 3 mosvc3_CDNS_7246542145921 $T=223775 183420 1 0 $X=222975 $Y=157800
X16 2 3 mosvc3_CDNS_7246542145921 $T=223775 185680 0 0 $X=222975 $Y=185250
X17 2 3 mosvc3_CDNS_7246542145921 $T=256775 183420 1 0 $X=255975 $Y=157800
X18 2 3 mosvc3_CDNS_7246542145921 $T=256775 185680 0 0 $X=255975 $Y=185250
X19 2 3 mosvc3_CDNS_7246542145921 $T=289775 183420 1 0 $X=288975 $Y=157800
X20 2 3 mosvc3_CDNS_7246542145921 $T=289775 185680 0 0 $X=288975 $Y=185250
X21 2 3 mosvc3_CDNS_7246542145921 $T=322775 183420 1 0 $X=321975 $Y=157800
X22 2 3 mosvc3_CDNS_7246542145921 $T=322775 185680 0 0 $X=321975 $Y=185250
X23 2 3 mosvc3_CDNS_7246542145921 $T=355775 183420 1 0 $X=354975 $Y=157800
X24 2 3 mosvc3_CDNS_7246542145921 $T=355775 185680 0 0 $X=354975 $Y=185250
X25 2 3 mosvc3_CDNS_7246542145921 $T=388775 183420 1 0 $X=387975 $Y=157800
X26 2 3 mosvc3_CDNS_7246542145921 $T=388775 185680 0 0 $X=387975 $Y=185250
X27 2 3 mosvc3_CDNS_7246542145921 $T=421775 183420 1 0 $X=420975 $Y=157800
X28 2 3 mosvc3_CDNS_7246542145921 $T=421775 185680 0 0 $X=420975 $Y=185250
X29 2 3 1 8 9 constant_gm $T=6360 5750 0 0 $X=7225 $Y=6590
.ends bias
