* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : pulse_generator                              *
* Netlisted  : Mon Aug 26 08:47:03 2024                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 LDDN(nedia) nedia2_d dnwtrm(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 1 MN(ne3) nem ndiff(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 2 MP(pe3) pem pdiff(D) p1trm(G) pdiff(S) nwtrm(B)
*.DEVTMPLT 3 NE3I_6() nemi_6 ndiff(D) p1trm(G) ndiff(S) pwitrm(B) dnwtrm(NW) bulk(SB)
*.DEVTMPLT 4 MOSVC3() mosvcm p1trm(G) nwtrm(NW) bulk(SB)
*.DEVTMPLT 5 R(s_res) s_res bulk(POS) bulk(NEG)
*.DEVTMPLT 6 D(p_dnw) p_dnw bulk(POS) nwtrm(NEG)
*.DEVTMPLT 7 D(p_ddnw) p_ddnw bulk(POS) dnwtrm(NEG)
*.DEVTMPLT 8 D(p_dipdnwmv) p_dipwmv pwitrm(POS) dnwtrm(NEG)
*.DEVTMPLT 9 D(p_dnw3) p_dnwm bulk(POS) nwtrm(NEG)
*.DEVTMPLT 10 R(rpp1k1_3) rpp1k1_s p1trm(POS) p1trm(NEG) bulk(SUB)
*.DEVTMPLT 11 R(rpp1k1_3) rpp1k1_n p1trm(POS) p1trm(NEG) nwtrm(SUB)
*.DEVTMPLT 12 C(cmm5t) cmim capm(POS) m4trm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NE3I_6                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NE3I_6 D G S B NW SB
.ends NE3I_6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MOSVC3                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MOSVC3 G NW SB
.ends MOSVC3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: LDDN                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt LDDN D G S B
.ends LDDN

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724654816050                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724654816050 1 2 3
** N=3 EP=3 FDC=4
M0 3 2 1 1 ne3 L=5e-07 W=5e-06 AD=1.35e-12 AS=2.4e-12 PD=5.54e-06 PS=1.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 1 ne3 L=5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=1040 $Y=0 $dt=1
M2 3 2 1 1 ne3 L=5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=2080 $Y=0 $dt=1
M3 1 2 3 1 ne3 L=5e-07 W=5e-06 AD=2.4e-12 AS=1.35e-12 PD=1.096e-05 PS=5.54e-06 $X=3120 $Y=0 $dt=1
.ends ne3_CDNS_724654816050

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nedia_CDNS_724654816051                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nedia_CDNS_724654816051 1 2 3 4
** N=4 EP=4 FDC=1
X0 2 4 3 1 LDDN w=5e-05 l=1.25e-06 adio=1.08602e-09 pdio=0.00013535 extlay=1 $[nedia] $X=-680 $Y=-4850 $dt=0
.ends nedia_CDNS_724654816051

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724654816052                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724654816052 1 2 3
** N=3 EP=3 FDC=4
M0 3 2 1 1 ne3 L=3.5e-07 W=5e-06 AD=1.35e-12 AS=2.4e-12 PD=5.54e-06 PS=1.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 1 ne3 L=3.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=890 $Y=0 $dt=1
M2 3 2 1 1 ne3 L=3.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=1780 $Y=0 $dt=1
M3 1 2 3 1 ne3 L=3.5e-07 W=5e-06 AD=2.4e-12 AS=1.35e-12 PD=1.096e-05 PS=5.54e-06 $X=2670 $Y=0 $dt=1
.ends ne3_CDNS_724654816052

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_724654816053                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_724654816053 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.00010265 W=4e-06 $[rpp1k1_3] $SUB=3 $X=0 $Y=0 $dt=10
.ends rpp1k1_3_CDNS_724654816053

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nedia_CDNS_724654816054                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nedia_CDNS_724654816054 1 2 3 4
** N=4 EP=4 FDC=8
X0 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=-680 $Y=-4850 $dt=0
X1 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=11220 $Y=-4850 $dt=0
X2 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=23120 $Y=-4850 $dt=0
X3 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=35020 $Y=-4850 $dt=0
X4 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=46920 $Y=-4850 $dt=0
X5 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=58820 $Y=-4850 $dt=0
X6 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=70720 $Y=-4850 $dt=0
X7 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=82620 $Y=-4850 $dt=0
.ends nedia_CDNS_724654816054

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724654816055                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724654816055 1 2 3 4
** N=4 EP=4 FDC=2
M0 3 2 1 4 ne3 L=1e-05 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 ne3 L=1e-05 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=10540 $Y=0 $dt=1
.ends ne3_CDNS_724654816055

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724654816056                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724654816056 1 2 3 4
*.DEVICECLIMB
** N=5 EP=4 FDC=1
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
.ends pe3_CDNS_724654816056

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724654816057                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724654816057 1 2 3
*.DEVICECLIMB
** N=4 EP=3 FDC=2
M0 3 2 1 1 pe3 L=3e-07 W=3e-06 AD=8.1e-13 AS=1.44e-12 PD=3.54e-06 PS=6.96e-06 $X=0 $Y=0 $dt=2
M1 1 2 3 1 pe3 L=3e-07 W=3e-06 AD=1.44e-12 AS=8.1e-13 PD=6.96e-06 PS=3.54e-06 $X=840 $Y=0 $dt=2
.ends pe3_CDNS_724654816057

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_724654816058                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_724654816058 1 2 3
** N=3 EP=3 FDC=1
R0 1 2 L=0.00204354 W=2e-06 $[rpp1k1_3] $SUB=3 $X=-2220 $Y=0 $dt=10
.ends rpp1k1_3_CDNS_724654816058

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160511                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160511 1 2 3 4
*.DEVICECLIMB
** N=5 EP=4 FDC=1
M0 3 2 1 4 pe3 L=5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
.ends pe3_CDNS_7246548160511

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7246548160512                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7246548160512 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=1e-05 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends ne3_CDNS_7246548160512

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7246548160513                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7246548160513 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=1e-06 W=5e-06 AD=2.4e-12 AS=2.4e-12 PD=1.096e-05 PS=1.096e-05 $X=0 $Y=0 $dt=1
.ends ne3_CDNS_7246548160513

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160514                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160514 1 2 3
*.DEVICECLIMB
** N=3 EP=3 FDC=9
M0 3 2 1 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
M1 1 2 3 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=5540 $Y=0 $dt=2
M2 3 2 1 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=11080 $Y=0 $dt=2
M3 1 2 3 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=16620 $Y=0 $dt=2
M4 3 2 1 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=22160 $Y=0 $dt=2
M5 1 2 3 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=27700 $Y=0 $dt=2
M6 3 2 1 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=33240 $Y=0 $dt=2
M7 1 2 3 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=38780 $Y=0 $dt=2
M8 3 2 1 1 pe3 L=5e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=44320 $Y=0 $dt=2
.ends pe3_CDNS_7246548160514

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7246548160515                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7246548160515 1 2 3
** N=3 EP=3 FDC=1
R0 1 2 L=1e-05 W=2e-06 $[rpp1k1_3] $SUB=3 $X=0 $Y=0 $dt=10
.ends rpp1k1_3_CDNS_7246548160515

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7246548160516                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7246548160516 1 2 3
*.DEVICECLIMB
** N=4 EP=3 FDC=1
R0 2 1 L=0.00016435 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=11
.ends rpp1k1_3_CDNS_7246548160516

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7246548160517                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7246548160517 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.00041122 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=10
.ends rpp1k1_3_CDNS_7246548160517

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7246548160518                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7246548160518 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=3.5e-07 W=2e-06 AD=9.6e-13 AS=9.6e-13 PD=4.96e-06 PS=4.96e-06 $X=0 $Y=0 $dt=1
.ends ne3_CDNS_7246548160518

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: current_source_gm_10_en_r                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt current_source_gm_10_en_r GNDA VDD3A EN BIAS PACTIVE IN FB VSUBHV GNDHV VDDHV
+ OUT
*.DEVICECLIMB
** N=27 EP=11 FDC=197
X404 GNDA 20 19 ne3_CDNS_724654816050 $T=248120 21400 0 0 $X=247320 $Y=21000
X405 VSUBHV 23 GNDHV 19 nedia_CDNS_724654816051 $T=282450 37820 0 0 $X=266230 $Y=18430
X406 GNDA 26 12 ne3_CDNS_724654816052 $T=25060 81535 0 0 $X=24260 $Y=80955
X407 GNDA 25 20 ne3_CDNS_724654816052 $T=30635 81535 0 0 $X=29835 $Y=80955
X408 23 GNDHV VSUBHV rpp1k1_3_CDNS_724654816053 $T=317545 27490 0 90 $X=309065 $Y=26550
X409 VSUBHV OUT FB 23 nedia_CDNS_724654816054 $T=441980 141045 0 270 $X=422590 $Y=41525
X410 12 BIAS BIAS GNDA ne3_CDNS_724654816055 $T=8060 64240 0 0 $X=7260 $Y=63840
X411 13 BIAS 14 GNDA ne3_CDNS_724654816055 $T=33845 64240 0 0 $X=33045 $Y=63840
X412 15 BIAS 16 GNDA ne3_CDNS_724654816055 $T=59570 64240 0 0 $X=58770 $Y=63840
X413 VDD3A 14 19 VDD3A pe3_CDNS_724654816056 $T=63965 94930 0 180 $X=61455 $Y=83900
X414 VDD3A 14 19 VDD3A pe3_CDNS_724654816056 $T=66205 94930 0 180 $X=63695 $Y=83900
X415 VDD3A 14 14 VDD3A pe3_CDNS_724654816056 $T=68445 94930 0 180 $X=65935 $Y=83900
X416 VDD3A 14 19 VDD3A pe3_CDNS_724654816056 $T=70685 94930 0 180 $X=68175 $Y=83900
X417 VDD3A 14 19 VDD3A pe3_CDNS_724654816056 $T=72925 94930 0 180 $X=70415 $Y=83900
X418 VDD3A EN 26 pe3_CDNS_724654816057 $T=15530 89865 0 180 $X=13480 $Y=86295
X419 VDD3A PACTIVE 25 pe3_CDNS_724654816057 $T=19690 89865 0 180 $X=17640 $Y=86295
X420 GNDHV OUT VSUBHV rpp1k1_3_CDNS_724654816058 $T=558265 45130 0 90 $X=515365 $Y=41970
X421 VDD3A VDD3A VDD3A VDD3A pe3_CDNS_7246548160511 $T=109700 69700 0 0 $X=108190 $Y=68670
X422 VDD3A VDD3A VDD3A VDD3A pe3_CDNS_7246548160511 $T=109700 93320 1 0 $X=108190 $Y=82290
X423 VDD3A VDD3A VDD3A VDD3A pe3_CDNS_7246548160511 $T=113660 125985 0 0 $X=112150 $Y=124955
X424 VDD3A VDD3A VDD3A VDD3A pe3_CDNS_7246548160511 $T=113660 148965 1 0 $X=112150 $Y=137935
X425 22 18 20 VDD3A pe3_CDNS_7246548160511 $T=115940 69700 0 0 $X=114430 $Y=68670
X426 22 17 21 VDD3A pe3_CDNS_7246548160511 $T=115940 93320 1 0 $X=114430 $Y=82290
X427 VDD3A 16 22 VDD3A pe3_CDNS_7246548160511 $T=119900 125985 0 0 $X=118390 $Y=124955
X428 VDD3A 16 22 VDD3A pe3_CDNS_7246548160511 $T=119900 148965 1 0 $X=118390 $Y=137935
X429 22 17 21 VDD3A pe3_CDNS_7246548160511 $T=122180 69700 0 0 $X=120670 $Y=68670
X430 22 18 20 VDD3A pe3_CDNS_7246548160511 $T=122180 93320 1 0 $X=120670 $Y=82290
X431 VDD3A 16 22 VDD3A pe3_CDNS_7246548160511 $T=126140 125985 0 0 $X=124630 $Y=124955
X432 VDD3A 16 22 VDD3A pe3_CDNS_7246548160511 $T=126140 148965 1 0 $X=124630 $Y=137935
X433 22 18 20 VDD3A pe3_CDNS_7246548160511 $T=128420 69700 0 0 $X=126910 $Y=68670
X434 22 17 21 VDD3A pe3_CDNS_7246548160511 $T=128420 93320 1 0 $X=126910 $Y=82290
X435 VDD3A 16 22 VDD3A pe3_CDNS_7246548160511 $T=132380 125985 0 0 $X=130870 $Y=124955
X436 VDD3A 16 22 VDD3A pe3_CDNS_7246548160511 $T=132380 148965 1 0 $X=130870 $Y=137935
X437 22 17 21 VDD3A pe3_CDNS_7246548160511 $T=134660 69700 0 0 $X=133150 $Y=68670
X438 22 18 20 VDD3A pe3_CDNS_7246548160511 $T=134660 93320 1 0 $X=133150 $Y=82290
X439 VDD3A 16 22 VDD3A pe3_CDNS_7246548160511 $T=138620 125985 0 0 $X=137110 $Y=124955
X440 VDD3A 16 22 VDD3A pe3_CDNS_7246548160511 $T=138620 148965 1 0 $X=137110 $Y=137935
X441 22 18 20 VDD3A pe3_CDNS_7246548160511 $T=140900 69700 0 0 $X=139390 $Y=68670
X442 22 17 21 VDD3A pe3_CDNS_7246548160511 $T=140900 93320 1 0 $X=139390 $Y=82290
X443 VDD3A 16 22 VDD3A pe3_CDNS_7246548160511 $T=144860 125985 0 0 $X=143350 $Y=124955
X444 VDD3A 16 22 VDD3A pe3_CDNS_7246548160511 $T=144860 148965 1 0 $X=143350 $Y=137935
X445 22 17 21 VDD3A pe3_CDNS_7246548160511 $T=147140 69700 0 0 $X=145630 $Y=68670
X446 22 18 20 VDD3A pe3_CDNS_7246548160511 $T=147140 93320 1 0 $X=145630 $Y=82290
X447 VDD3A 16 18 VDD3A pe3_CDNS_7246548160511 $T=151100 125985 0 0 $X=149590 $Y=124955
X448 VDD3A 16 17 VDD3A pe3_CDNS_7246548160511 $T=151100 148965 1 0 $X=149590 $Y=137935
X449 22 18 20 VDD3A pe3_CDNS_7246548160511 $T=153380 69700 0 0 $X=151870 $Y=68670
X450 22 17 21 VDD3A pe3_CDNS_7246548160511 $T=153380 93320 1 0 $X=151870 $Y=82290
X451 VDD3A 16 16 VDD3A pe3_CDNS_7246548160511 $T=157340 125985 0 0 $X=155830 $Y=124955
X452 VDD3A 16 16 VDD3A pe3_CDNS_7246548160511 $T=157340 148965 1 0 $X=155830 $Y=137935
X453 22 17 21 VDD3A pe3_CDNS_7246548160511 $T=159620 69700 0 0 $X=158110 $Y=68670
X454 22 18 20 VDD3A pe3_CDNS_7246548160511 $T=159620 93320 1 0 $X=158110 $Y=82290
X455 VDD3A 16 17 VDD3A pe3_CDNS_7246548160511 $T=163580 125985 0 0 $X=162070 $Y=124955
X456 VDD3A 16 18 VDD3A pe3_CDNS_7246548160511 $T=163580 148965 1 0 $X=162070 $Y=137935
X457 22 18 20 VDD3A pe3_CDNS_7246548160511 $T=165860 69700 0 0 $X=164350 $Y=68670
X458 22 17 21 VDD3A pe3_CDNS_7246548160511 $T=165860 93320 1 0 $X=164350 $Y=82290
X459 VDD3A 16 22 VDD3A pe3_CDNS_7246548160511 $T=169820 125985 0 0 $X=168310 $Y=124955
X460 VDD3A 16 22 VDD3A pe3_CDNS_7246548160511 $T=169820 148965 1 0 $X=168310 $Y=137935
X461 22 17 21 VDD3A pe3_CDNS_7246548160511 $T=172100 69700 0 0 $X=170590 $Y=68670
X462 22 18 20 VDD3A pe3_CDNS_7246548160511 $T=172100 93320 1 0 $X=170590 $Y=82290
X463 VDD3A 16 22 VDD3A pe3_CDNS_7246548160511 $T=176060 125985 0 0 $X=174550 $Y=124955
X464 VDD3A 16 22 VDD3A pe3_CDNS_7246548160511 $T=176060 148965 1 0 $X=174550 $Y=137935
X465 22 18 20 VDD3A pe3_CDNS_7246548160511 $T=178340 69700 0 0 $X=176830 $Y=68670
X466 22 17 21 VDD3A pe3_CDNS_7246548160511 $T=178340 93320 1 0 $X=176830 $Y=82290
X467 VDD3A 16 22 VDD3A pe3_CDNS_7246548160511 $T=182300 125985 0 0 $X=180790 $Y=124955
X468 VDD3A 16 22 VDD3A pe3_CDNS_7246548160511 $T=182300 148965 1 0 $X=180790 $Y=137935
X469 22 17 21 VDD3A pe3_CDNS_7246548160511 $T=184580 69700 0 0 $X=183070 $Y=68670
X470 22 18 20 VDD3A pe3_CDNS_7246548160511 $T=184580 93320 1 0 $X=183070 $Y=82290
X471 VDD3A 16 22 VDD3A pe3_CDNS_7246548160511 $T=188540 125985 0 0 $X=187030 $Y=124955
X472 VDD3A 16 22 VDD3A pe3_CDNS_7246548160511 $T=188540 148965 1 0 $X=187030 $Y=137935
X473 22 18 20 VDD3A pe3_CDNS_7246548160511 $T=190820 69700 0 0 $X=189310 $Y=68670
X474 22 17 21 VDD3A pe3_CDNS_7246548160511 $T=190820 93320 1 0 $X=189310 $Y=82290
X475 VDD3A 16 22 VDD3A pe3_CDNS_7246548160511 $T=194780 125985 0 0 $X=193270 $Y=124955
X476 VDD3A 16 22 VDD3A pe3_CDNS_7246548160511 $T=194780 148965 1 0 $X=193270 $Y=137935
X477 22 17 21 VDD3A pe3_CDNS_7246548160511 $T=197060 69700 0 0 $X=195550 $Y=68670
X478 22 18 20 VDD3A pe3_CDNS_7246548160511 $T=197060 93320 1 0 $X=195550 $Y=82290
X479 VDD3A VDD3A VDD3A VDD3A pe3_CDNS_7246548160511 $T=201020 125985 0 0 $X=199510 $Y=124955
X480 VDD3A VDD3A VDD3A VDD3A pe3_CDNS_7246548160511 $T=201020 148965 1 0 $X=199510 $Y=137935
X481 VDD3A VDD3A VDD3A VDD3A pe3_CDNS_7246548160511 $T=203300 69700 0 0 $X=201790 $Y=68670
X482 VDD3A VDD3A VDD3A VDD3A pe3_CDNS_7246548160511 $T=203300 93320 1 0 $X=201790 $Y=82290
X483 GNDA GNDA GNDA ne3_CDNS_7246548160512 $T=17420 20740 0 0 $X=16620 $Y=20340
X484 GNDA GNDA GNDA ne3_CDNS_7246548160512 $T=17420 42860 1 0 $X=16620 $Y=32290
X485 GNDA 12 15 ne3_CDNS_7246548160512 $T=28660 20740 0 0 $X=27860 $Y=20340
X486 GNDA 12 15 ne3_CDNS_7246548160512 $T=28660 42860 1 0 $X=27860 $Y=32290
X487 GNDA 12 12 ne3_CDNS_7246548160512 $T=39900 20740 0 0 $X=39100 $Y=20340
X488 GNDA 12 12 ne3_CDNS_7246548160512 $T=39900 42860 1 0 $X=39100 $Y=32290
X489 GNDA 12 13 ne3_CDNS_7246548160512 $T=51140 20740 0 0 $X=50340 $Y=20340
X490 GNDA 12 13 ne3_CDNS_7246548160512 $T=51140 42860 1 0 $X=50340 $Y=32290
X491 GNDA GNDA GNDA ne3_CDNS_7246548160512 $T=62380 20740 0 0 $X=61580 $Y=20340
X492 GNDA GNDA GNDA ne3_CDNS_7246548160512 $T=62380 42860 1 0 $X=61580 $Y=32290
X493 GNDA 21 20 ne3_CDNS_7246548160513 $T=232175 21040 0 0 $X=231375 $Y=20640
X494 GNDA 21 21 ne3_CDNS_7246548160513 $T=232175 32430 1 0 $X=231375 $Y=26860
X495 GNDA 21 21 ne3_CDNS_7246548160513 $T=234415 21040 0 0 $X=233615 $Y=20640
X496 GNDA 21 20 ne3_CDNS_7246548160513 $T=234415 32430 1 0 $X=233615 $Y=26860
X497 17 IN GNDA pe3_CDNS_7246548160514 $T=106815 19890 0 0 $X=105305 $Y=18860
X498 18 24 GNDA pe3_CDNS_7246548160514 $T=106815 43890 1 0 $X=105305 $Y=32860
X499 18 24 GNDA pe3_CDNS_7246548160514 $T=161095 19890 0 0 $X=159585 $Y=18860
X500 17 IN GNDA pe3_CDNS_7246548160514 $T=161095 43890 1 0 $X=159585 $Y=32860
X501 FB 24 GNDA rpp1k1_3_CDNS_7246548160515 $T=229190 61300 0 90 $X=226970 $Y=60360
X502 FB 24 GNDA rpp1k1_3_CDNS_7246548160515 $T=232060 61300 0 90 $X=229840 $Y=60360
X503 FB 24 GNDA rpp1k1_3_CDNS_7246548160515 $T=234930 61300 0 90 $X=232710 $Y=60360
X504 FB 24 GNDA rpp1k1_3_CDNS_7246548160515 $T=237800 61300 0 90 $X=235580 $Y=60360
X505 FB 24 GNDA rpp1k1_3_CDNS_7246548160515 $T=240670 61300 0 90 $X=238450 $Y=60360
X506 FB 24 GNDA rpp1k1_3_CDNS_7246548160515 $T=243540 61300 0 90 $X=241320 $Y=60360
X507 FB 24 GNDA rpp1k1_3_CDNS_7246548160515 $T=246410 61300 0 90 $X=244190 $Y=60360
X508 FB 24 GNDA rpp1k1_3_CDNS_7246548160515 $T=249280 61300 0 90 $X=247060 $Y=60360
X509 FB 24 GNDA rpp1k1_3_CDNS_7246548160515 $T=252150 61300 0 90 $X=249930 $Y=60360
X510 19 27 VDD3A rpp1k1_3_CDNS_7246548160516 $T=255085 124550 0 180 $X=228430 $Y=99030
X511 VDDHV 23 VSUBHV rpp1k1_3_CDNS_7246548160517 $T=322885 76685 0 270 $X=322665 $Y=25845
X512 GNDA EN 26 ne3_CDNS_7246548160518 $T=14340 81020 0 0 $X=13540 $Y=80620
X513 GNDA PACTIVE 25 ne3_CDNS_7246548160518 $T=18500 81020 0 0 $X=17700 $Y=80620
X756 VDD3A GNDA GNDA MOSVC3 w=2e-05 l=3e-05 $X=16180 $Y=110530 $dt=4
X757 VDD3A GNDA GNDA MOSVC3 w=2e-05 l=3e-05 $X=16180 $Y=132530 $dt=4
X758 VDD3A GNDA GNDA MOSVC3 w=2e-05 l=3e-05 $X=48780 $Y=110530 $dt=4
X759 VDD3A GNDA GNDA MOSVC3 w=2e-05 l=3e-05 $X=48780 $Y=132530 $dt=4
D4 GNDA VDD3A p_dnw AREA=3.57048e-11 PJ=3.588e-05 perimeter=3.588e-05 $X=11740 $Y=84695 $dt=6
D5 GNDA VDD3A p_dnw AREA=1.90124e-10 PJ=7.516e-05 perimeter=7.516e-05 $X=59815 $Y=81480 $dt=6
D6 GNDA VDD3A p_dnw AREA=1.58288e-09 PJ=0.00049318 perimeter=0.00049318 $X=99710 $Y=59910 $dt=6
D7 GNDA VDD3A p_dnw AREA=3.09086e-09 PJ=0.00032604 perimeter=0.00032604 $X=101390 $Y=114415 $dt=6
D8 GNDA 17 p_dnw AREA=1.82058e-10 PJ=5.826e-05 perimeter=5.826e-05 $X=105905 $Y=15300 $dt=6
D9 GNDA 18 p_dnw AREA=1.82058e-10 PJ=5.826e-05 perimeter=5.826e-05 $X=105905 $Y=44920 $dt=6
D10 GNDA 18 p_dnw AREA=1.82058e-10 PJ=5.826e-05 perimeter=5.826e-05 $X=160185 $Y=15300 $dt=6
D11 GNDA 17 p_dnw AREA=1.82058e-10 PJ=5.826e-05 perimeter=5.826e-05 $X=160185 $Y=44920 $dt=6
D12 GNDA VDD3A p_dnw AREA=8.36476e-09 PJ=0.0003905 perimeter=0.0003905 $X=226790 $Y=95600 $dt=6
D13 GNDA VDD3A p_dnw3 AREA=4.20992e-11 PJ=0 perimeter=0 $X=12880 $Y=85835 $dt=9
D14 GNDA GNDA p_dnw3 AREA=5.9176e-11 PJ=0.00010492 perimeter=0.00010492 $X=15380 $Y=110100 $dt=9
D15 GNDA GNDA p_dnw3 AREA=5.9176e-11 PJ=0.00010492 perimeter=0.00010492 $X=15380 $Y=132100 $dt=9
D16 GNDA GNDA p_dnw3 AREA=5.9176e-11 PJ=0.00010492 perimeter=0.00010492 $X=47980 $Y=110100 $dt=9
D17 GNDA GNDA p_dnw3 AREA=5.9176e-11 PJ=0.00010492 perimeter=0.00010492 $X=47980 $Y=132100 $dt=9
D18 GNDA VDD3A p_dnw3 AREA=1.56539e-10 PJ=0 perimeter=0 $X=61455 $Y=83900 $dt=9
D19 GNDA 17 p_dnw3 AREA=5.86064e-10 PJ=7.406e-05 perimeter=7.406e-05 $X=105905 $Y=18860 $dt=9
D20 GNDA 18 p_dnw3 AREA=5.86064e-10 PJ=7.406e-05 perimeter=7.406e-05 $X=105905 $Y=33460 $dt=9
D21 GNDA VDD3A p_dnw3 AREA=1.22554e-09 PJ=0 perimeter=0 $X=108190 $Y=68670 $dt=9
D22 GNDA VDD3A p_dnw3 AREA=1.15225e-09 PJ=0.00012214 perimeter=0.00012214 $X=108190 $Y=82290 $dt=9
D23 GNDA VDD3A p_dnw3 AREA=1.15028e-09 PJ=0 perimeter=0 $X=112150 $Y=124955 $dt=9
D24 GNDA VDD3A p_dnw3 AREA=1.15028e-09 PJ=0 perimeter=0 $X=112150 $Y=137935 $dt=9
D25 GNDA 18 p_dnw3 AREA=5.86064e-10 PJ=7.406e-05 perimeter=7.406e-05 $X=160185 $Y=18860 $dt=9
D26 GNDA 17 p_dnw3 AREA=5.86064e-10 PJ=7.406e-05 perimeter=7.406e-05 $X=160185 $Y=33460 $dt=9
C27 20 27 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=231620 $Y=128940 $dt=12
C28 20 27 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=263220 $Y=97740 $dt=12
C29 20 27 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=263220 $Y=128940 $dt=12
C30 20 27 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=294820 $Y=97740 $dt=12
C31 20 27 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=294820 $Y=128940 $dt=12
C32 20 27 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=326420 $Y=97740 $dt=12
C33 20 27 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=326420 $Y=128940 $dt=12
.ends current_source_gm_10_en_r

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: mosvc3_CDNS_7246548160521                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt mosvc3_CDNS_7246548160521 1 2
** N=2 EP=2 FDC=2
X0 2 1 1 MOSVC3 w=2.5e-05 l=2e-05 $X=0 $Y=0 $dt=4
D1 1 1 p_dnw3 AREA=5.8576e-11 PJ=9.492e-05 perimeter=9.492e-05 $X=-800 $Y=-430 $dt=9
.ends mosvc3_CDNS_7246548160521

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: mosvc3_CDNS_7246548160522                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt mosvc3_CDNS_7246548160522 1 2
** N=2 EP=2 FDC=2
X0 2 1 1 MOSVC3 w=2e-05 l=2e-05 $X=0 $Y=0 $dt=4
D1 1 1 p_dnw3 AREA=5.0576e-11 PJ=8.492e-05 perimeter=8.492e-05 $X=-800 $Y=-430 $dt=9
.ends mosvc3_CDNS_7246548160522

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160523                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160523 1 2 3
*.DEVICECLIMB
** N=4 EP=3 FDC=1
M0 3 2 1 1 pe3 L=1e-05 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
.ends pe3_CDNS_7246548160523

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160524                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160524 1 2 3 4
*.DEVICECLIMB
** N=5 EP=4 FDC=2
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=2
.ends pe3_CDNS_7246548160524

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160525                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160525 1 2 3 4
*.DEVICECLIMB
** N=5 EP=4 FDC=4
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=2
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=2
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=2
.ends pe3_CDNS_7246548160525

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160526                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160526 1 2 3 4
*.DEVICECLIMB
** N=5 EP=4 FDC=8
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=2
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=2
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=2
M4 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=6160 $Y=0 $dt=2
M5 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7700 $Y=0 $dt=2
M6 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=9240 $Y=0 $dt=2
M7 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=10780 $Y=0 $dt=2
.ends pe3_CDNS_7246548160526

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160527                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160527 1 2 3 4
*.DEVICECLIMB
** N=5 EP=4 FDC=16
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=2
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=2
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=2
M4 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=6160 $Y=0 $dt=2
M5 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7700 $Y=0 $dt=2
M6 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=9240 $Y=0 $dt=2
M7 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10780 $Y=0 $dt=2
M8 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12320 $Y=0 $dt=2
M9 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=13860 $Y=0 $dt=2
M10 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=15400 $Y=0 $dt=2
M11 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=16940 $Y=0 $dt=2
M12 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=18480 $Y=0 $dt=2
M13 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=20020 $Y=0 $dt=2
M14 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=21560 $Y=0 $dt=2
M15 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=23100 $Y=0 $dt=2
.ends pe3_CDNS_7246548160527

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160528                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160528 1 2 3 4
*.DEVICECLIMB
** N=5 EP=4 FDC=32
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=2
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=2
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=2
M4 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=6160 $Y=0 $dt=2
M5 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7700 $Y=0 $dt=2
M6 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=9240 $Y=0 $dt=2
M7 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10780 $Y=0 $dt=2
M8 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12320 $Y=0 $dt=2
M9 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=13860 $Y=0 $dt=2
M10 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=15400 $Y=0 $dt=2
M11 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=16940 $Y=0 $dt=2
M12 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=18480 $Y=0 $dt=2
M13 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=20020 $Y=0 $dt=2
M14 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=21560 $Y=0 $dt=2
M15 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=23100 $Y=0 $dt=2
M16 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=24640 $Y=0 $dt=2
M17 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=26180 $Y=0 $dt=2
M18 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=27720 $Y=0 $dt=2
M19 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=29260 $Y=0 $dt=2
M20 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=30800 $Y=0 $dt=2
M21 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=32340 $Y=0 $dt=2
M22 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=33880 $Y=0 $dt=2
M23 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=35420 $Y=0 $dt=2
M24 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=36960 $Y=0 $dt=2
M25 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=38500 $Y=0 $dt=2
M26 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=40040 $Y=0 $dt=2
M27 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=41580 $Y=0 $dt=2
M28 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=43120 $Y=0 $dt=2
M29 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=44660 $Y=0 $dt=2
M30 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=46200 $Y=0 $dt=2
M31 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=47740 $Y=0 $dt=2
.ends pe3_CDNS_7246548160528

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7246548160529                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7246548160529 1 2
** N=2 EP=2 FDC=1
R0 2 1 L=0.00021702 W=4e-06 $[rpp1k1_3] $SUB=2 $X=-4220 $Y=0 $dt=10
.ends rpp1k1_3_CDNS_7246548160529

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160530                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160530 1 2 3 4
*.DEVICECLIMB
** N=5 EP=4 FDC=10
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=2
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=2
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=2
M4 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=6160 $Y=0 $dt=2
M5 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7700 $Y=0 $dt=2
M6 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=9240 $Y=0 $dt=2
M7 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10780 $Y=0 $dt=2
M8 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12320 $Y=0 $dt=2
M9 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=13860 $Y=0 $dt=2
.ends pe3_CDNS_7246548160530

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7246548160531                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7246548160531 1 2
** N=2 EP=2 FDC=1
R0 2 1 L=0.0008227 W=4e-06 $[rpp1k1_3] $SUB=2 $X=-4220 $Y=0 $dt=10
.ends rpp1k1_3_CDNS_7246548160531

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160532                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160532 1 2
*.DEVICECLIMB
** N=3 EP=2 FDC=1
M0 2 2 1 1 pe3 L=2e-05 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
.ends pe3_CDNS_7246548160532

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160533                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160533 1 2 3
*.DEVICECLIMB
** N=4 EP=3 FDC=1
M0 3 2 1 1 pe3 L=3e-07 W=6e-06 AD=2.88e-12 AS=2.88e-12 PD=1.296e-05 PS=1.296e-05 $X=0 $Y=0 $dt=2
.ends pe3_CDNS_7246548160533

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160534                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160534 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=2
M0 3 2 1 4 pe3 L=3.5e-07 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
M1 1 2 3 4 pe3 L=3.5e-07 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=890 $Y=0 $dt=2
.ends pe3_CDNS_7246548160534

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7246548160535                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7246548160535 1 2 3 4
** N=4 EP=4 FDC=8
M0 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=2540 $Y=0 $dt=1
M2 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=5080 $Y=0 $dt=1
M3 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7620 $Y=0 $dt=1
M4 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10160 $Y=0 $dt=1
M5 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12700 $Y=0 $dt=1
M6 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=15240 $Y=0 $dt=1
M7 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=17780 $Y=0 $dt=1
.ends ne3_CDNS_7246548160535

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3i_6_CDNS_7246548160536                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3i_6_CDNS_7246548160536 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=1
X0 1 2 3 1 4 5 NE3I_6 w=1e-05 l=2e-06 as=4.8e-12 ad=4.8e-12 ps=2.096e-05 pd=2.096e-05 $X=0 $Y=0 $dt=3
.ends ne3i_6_CDNS_7246548160536

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7246548160537                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7246548160537 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=2e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends ne3_CDNS_7246548160537

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160538                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160538 1
*.DEVICECLIMB
** N=2 EP=1 FDC=1
M0 1 1 1 1 pe3 L=1e-05 W=2e-06 AD=9.6e-13 AS=9.6e-13 PD=4.96e-06 PS=4.96e-06 $X=0 $Y=0 $dt=2
.ends pe3_CDNS_7246548160538

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7246548160539                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7246548160539 1 2 3
** N=3 EP=3 FDC=4
M0 3 2 1 1 ne3 L=3.5e-07 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 1 ne3 L=3.5e-07 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=890 $Y=0 $dt=1
M2 3 2 1 1 ne3 L=3.5e-07 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1780 $Y=0 $dt=1
M3 1 2 3 1 ne3 L=3.5e-07 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=2670 $Y=0 $dt=1
.ends ne3_CDNS_7246548160539

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A15                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A15 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=8 EP=7 FDC=4
X0 3 2 1 pe3_CDNS_7246548160523 $T=1510 11030 1 0 $X=0 $Y=0
X1 3 5 4 pe3_CDNS_7246548160523 $T=12750 11030 1 0 $X=11240 $Y=0
X2 3 5 6 pe3_CDNS_7246548160523 $T=23990 11030 1 0 $X=22480 $Y=0
X3 3 5 7 pe3_CDNS_7246548160523 $T=35230 11030 1 0 $X=33720 $Y=0
.ends MASCO__A15

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: dac6b_amp_n2                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt dac6b_amp_n2 GNDA VDDA BIAS ENABLE VOUT VREF D5 D4 D3 D2
+ D1 D0
** N=31 EP=12 FDC=372
X280 24 19 VOUT VDDA pe3_CDNS_724654816056 $T=373510 36320 1 0 $X=372000 $Y=25290
X281 GNDA ENABLE 25 ne3_CDNS_7246548160518 $T=91035 56560 0 0 $X=90235 $Y=56160
X1107 VDDA 15 15 pe3_CDNS_7246548160523 $T=15710 148580 0 0 $X=14200 $Y=147550
X1108 VDDA 15 20 pe3_CDNS_7246548160523 $T=15710 171560 1 0 $X=14200 $Y=160530
X1109 VDDA 15 20 pe3_CDNS_7246548160523 $T=26950 148580 0 0 $X=25440 $Y=147550
X1110 VDDA 15 15 pe3_CDNS_7246548160523 $T=26950 171560 1 0 $X=25440 $Y=160530
X1111 VDDA VDDA VDDA pe3_CDNS_7246548160523 $T=56340 148580 0 0 $X=54830 $Y=147550
X1112 VDDA 16 16 pe3_CDNS_7246548160523 $T=67580 148580 0 0 $X=66070 $Y=147550
X1113 VDDA 16 17 pe3_CDNS_7246548160523 $T=78820 148580 0 0 $X=77310 $Y=147550
X1114 VDDA 16 16 pe3_CDNS_7246548160523 $T=90060 148580 0 0 $X=88550 $Y=147550
X1115 VDDA 16 17 pe3_CDNS_7246548160523 $T=101300 148580 0 0 $X=99790 $Y=147550
X1116 VDDA 16 16 pe3_CDNS_7246548160523 $T=112540 148580 0 0 $X=111030 $Y=147550
X1117 VDDA 16 17 pe3_CDNS_7246548160523 $T=123780 148580 0 0 $X=122270 $Y=147550
X1118 VDDA 16 16 pe3_CDNS_7246548160523 $T=135020 148580 0 0 $X=133510 $Y=147550
X1119 VDDA 16 17 pe3_CDNS_7246548160523 $T=146260 148580 0 0 $X=144750 $Y=147550
X1120 VDDA 16 16 pe3_CDNS_7246548160523 $T=146260 171560 1 0 $X=144750 $Y=160530
X1121 VDDA VDDA VDDA pe3_CDNS_7246548160523 $T=157500 148580 0 0 $X=155990 $Y=147550
X1122 VDDA VDDA VDDA pe3_CDNS_7246548160523 $T=157500 171560 1 0 $X=155990 $Y=160530
X1123 VDDA VDDA VDDA pe3_CDNS_7246548160523 $T=340315 71115 1 0 $X=338805 $Y=60085
X1124 VDDA 17 26 pe3_CDNS_7246548160523 $T=340315 89915 1 0 $X=338805 $Y=78885
X1125 VDDA 17 26 pe3_CDNS_7246548160523 $T=340315 108715 1 0 $X=338805 $Y=97685
X1126 VDDA 17 26 pe3_CDNS_7246548160523 $T=340315 127515 1 0 $X=338805 $Y=116485
X1127 VDDA 17 26 pe3_CDNS_7246548160523 $T=340315 146315 1 0 $X=338805 $Y=135285
X1128 VDDA 17 26 pe3_CDNS_7246548160523 $T=340315 165115 1 0 $X=338805 $Y=154085
X1129 VDDA VDDA VDDA pe3_CDNS_7246548160523 $T=351555 71115 1 0 $X=350045 $Y=60085
X1130 VDDA 17 26 pe3_CDNS_7246548160523 $T=351555 89915 1 0 $X=350045 $Y=78885
X1131 VDDA 17 26 pe3_CDNS_7246548160523 $T=351555 108715 1 0 $X=350045 $Y=97685
X1132 VDDA 17 26 pe3_CDNS_7246548160523 $T=351555 127515 1 0 $X=350045 $Y=116485
X1133 VDDA 17 26 pe3_CDNS_7246548160523 $T=351555 146315 1 0 $X=350045 $Y=135285
X1134 VDDA 17 26 pe3_CDNS_7246548160523 $T=351555 165115 1 0 $X=350045 $Y=154085
X1135 VDDA VDDA VDDA pe3_CDNS_7246548160523 $T=362795 71115 1 0 $X=361285 $Y=60085
X1136 VDDA VDDA VDDA pe3_CDNS_7246548160523 $T=362795 89915 1 0 $X=361285 $Y=78885
X1137 VDDA VDDA VDDA pe3_CDNS_7246548160523 $T=362795 108715 1 0 $X=361285 $Y=97685
X1138 VDDA VDDA VDDA pe3_CDNS_7246548160523 $T=362795 127515 1 0 $X=361285 $Y=116485
X1139 VDDA VDDA VDDA pe3_CDNS_7246548160523 $T=362795 146315 1 0 $X=361285 $Y=135285
X1140 VDDA VDDA VDDA pe3_CDNS_7246548160523 $T=362795 165115 1 0 $X=361285 $Y=154085
X1141 29 19 VOUT VDDA pe3_CDNS_7246548160524 $T=364135 36320 1 0 $X=362625 $Y=25290
X1142 31 19 VOUT VDDA pe3_CDNS_7246548160525 $T=351800 36320 1 0 $X=350290 $Y=25290
X1143 28 19 VOUT VDDA pe3_CDNS_7246548160526 $T=333335 36320 1 0 $X=331825 $Y=25290
X1144 27 19 VOUT VDDA pe3_CDNS_7246548160527 $T=302570 36320 1 0 $X=301060 $Y=25290
X1145 26 19 VOUT VDDA pe3_CDNS_7246548160528 $T=246755 36320 1 0 $X=245245 $Y=25290
X1146 VOUT GNDA rpp1k1_3_CDNS_7246548160529 $T=190390 9160 0 0 $X=185230 $Y=8940
X1147 30 19 23 VDDA pe3_CDNS_7246548160530 $T=223935 36320 1 0 $X=222425 $Y=25290
X1148 23 GNDA rpp1k1_3_CDNS_7246548160531 $T=80195 9200 0 0 $X=75035 $Y=8980
X1149 18 GNDA pe3_CDNS_7246548160532 $T=154675 76695 0 0 $X=153165 $Y=75665
X1150 19 18 pe3_CDNS_7246548160532 $T=154675 98175 0 0 $X=153165 $Y=97145
X1151 20 19 pe3_CDNS_7246548160532 $T=154675 119125 0 0 $X=153165 $Y=118095
X1152 VDDA ENABLE 25 pe3_CDNS_7246548160533 $T=91085 67915 1 0 $X=90175 $Y=61345
X1153 26 D5 GNDA VDDA pe3_CDNS_7246548160534 $T=307075 17335 1 0 $X=305565 $Y=6305
X1154 27 D4 GNDA VDDA pe3_CDNS_7246548160534 $T=316335 17335 1 0 $X=314825 $Y=6305
X1155 28 D3 GNDA VDDA pe3_CDNS_7246548160534 $T=325595 17335 1 0 $X=324085 $Y=6305
X1156 31 D2 GNDA VDDA pe3_CDNS_7246548160534 $T=334855 17335 1 0 $X=333345 $Y=6305
X1157 29 D1 GNDA VDDA pe3_CDNS_7246548160534 $T=344115 17335 1 0 $X=342605 $Y=6305
X1158 24 D0 GNDA VDDA pe3_CDNS_7246548160534 $T=353375 17335 1 0 $X=351865 $Y=6305
X1159 13 BIAS BIAS GNDA ne3_CDNS_7246548160535 $T=7715 59435 0 0 $X=6915 $Y=59035
X1160 14 BIAS 15 GNDA ne3_CDNS_7246548160535 $T=34470 59435 0 0 $X=33670 $Y=59035
X1161 21 BIAS 22 GNDA ne3_CDNS_7246548160535 $T=62205 59435 0 0 $X=61405 $Y=59035
X1162 22 22 22 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=70370 100985 0 0 $X=66310 $Y=96535
X1163 22 22 22 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=70370 124285 1 0 $X=66310 $Y=109715
X1164 22 23 16 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=73770 100985 0 0 $X=69710 $Y=96535
X1165 22 VREF 17 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=73770 124285 1 0 $X=69710 $Y=109715
X1166 22 VREF 17 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=77170 100985 0 0 $X=73110 $Y=96535
X1167 22 23 16 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=77170 124285 1 0 $X=73110 $Y=109715
X1168 22 23 16 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=80570 100985 0 0 $X=76510 $Y=96535
X1169 22 VREF 17 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=80570 124285 1 0 $X=76510 $Y=109715
X1170 22 VREF 17 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=83970 100985 0 0 $X=79910 $Y=96535
X1171 22 23 16 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=83970 124285 1 0 $X=79910 $Y=109715
X1172 22 23 16 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=87370 100985 0 0 $X=83310 $Y=96535
X1173 22 VREF 17 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=87370 124285 1 0 $X=83310 $Y=109715
X1174 22 VREF 17 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=90770 100985 0 0 $X=86710 $Y=96535
X1175 22 23 16 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=90770 124285 1 0 $X=86710 $Y=109715
X1176 22 23 16 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=94170 100985 0 0 $X=90110 $Y=96535
X1177 22 VREF 17 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=94170 124285 1 0 $X=90110 $Y=109715
X1178 22 VREF 17 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=97570 100985 0 0 $X=93510 $Y=96535
X1179 22 23 16 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=97570 124285 1 0 $X=93510 $Y=109715
X1180 22 23 16 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=100970 100985 0 0 $X=96910 $Y=96535
X1181 22 VREF 17 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=100970 124285 1 0 $X=96910 $Y=109715
X1182 22 VREF 17 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=104370 100985 0 0 $X=100310 $Y=96535
X1183 22 23 16 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=104370 124285 1 0 $X=100310 $Y=109715
X1184 22 23 16 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=107770 100985 0 0 $X=103710 $Y=96535
X1185 22 VREF 17 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=107770 124285 1 0 $X=103710 $Y=109715
X1186 22 VREF 17 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=111170 100985 0 0 $X=107110 $Y=96535
X1187 22 23 16 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=111170 124285 1 0 $X=107110 $Y=109715
X1188 22 23 16 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=114570 100985 0 0 $X=110510 $Y=96535
X1189 22 VREF 17 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=114570 124285 1 0 $X=110510 $Y=109715
X1190 22 VREF 17 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=117970 100985 0 0 $X=113910 $Y=96535
X1191 22 23 16 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=117970 124285 1 0 $X=113910 $Y=109715
X1192 22 23 16 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=121370 100985 0 0 $X=117310 $Y=96535
X1193 22 VREF 17 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=121370 124285 1 0 $X=117310 $Y=109715
X1194 22 VREF 17 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=124770 100985 0 0 $X=120710 $Y=96535
X1195 22 23 16 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=124770 124285 1 0 $X=120710 $Y=109715
X1196 22 22 22 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=128170 100985 0 0 $X=124110 $Y=96535
X1197 22 22 22 VDDA GNDA ne3i_6_CDNS_7246548160536 $T=128170 124285 1 0 $X=124110 $Y=109715
X1198 GNDA GNDA GNDA ne3_CDNS_7246548160537 $T=11530 16320 0 0 $X=10730 $Y=15920
X1199 GNDA GNDA GNDA ne3_CDNS_7246548160537 $T=11530 38460 1 0 $X=10730 $Y=27890
X1200 GNDA 13 21 ne3_CDNS_7246548160537 $T=14770 16320 0 0 $X=13970 $Y=15920
X1201 GNDA 13 13 ne3_CDNS_7246548160537 $T=14770 38460 1 0 $X=13970 $Y=27890
X1202 GNDA 13 14 ne3_CDNS_7246548160537 $T=18010 16320 0 0 $X=17210 $Y=15920
X1203 GNDA 13 21 ne3_CDNS_7246548160537 $T=18010 38460 1 0 $X=17210 $Y=27890
X1204 GNDA 13 13 ne3_CDNS_7246548160537 $T=21250 16320 0 0 $X=20450 $Y=15920
X1205 GNDA 13 14 ne3_CDNS_7246548160537 $T=21250 38460 1 0 $X=20450 $Y=27890
X1206 GNDA 13 21 ne3_CDNS_7246548160537 $T=24490 16320 0 0 $X=23690 $Y=15920
X1207 GNDA 13 13 ne3_CDNS_7246548160537 $T=24490 38460 1 0 $X=23690 $Y=27890
X1208 GNDA 13 14 ne3_CDNS_7246548160537 $T=27730 16320 0 0 $X=26930 $Y=15920
X1209 GNDA 13 21 ne3_CDNS_7246548160537 $T=27730 38460 1 0 $X=26930 $Y=27890
X1210 GNDA 13 13 ne3_CDNS_7246548160537 $T=30970 16320 0 0 $X=30170 $Y=15920
X1211 GNDA 13 14 ne3_CDNS_7246548160537 $T=30970 38460 1 0 $X=30170 $Y=27890
X1212 GNDA 13 21 ne3_CDNS_7246548160537 $T=34210 16320 0 0 $X=33410 $Y=15920
X1213 GNDA 13 13 ne3_CDNS_7246548160537 $T=34210 38460 1 0 $X=33410 $Y=27890
X1214 GNDA 13 14 ne3_CDNS_7246548160537 $T=37450 16320 0 0 $X=36650 $Y=15920
X1215 GNDA 13 21 ne3_CDNS_7246548160537 $T=37450 38460 1 0 $X=36650 $Y=27890
X1216 GNDA 13 13 ne3_CDNS_7246548160537 $T=40690 16320 0 0 $X=39890 $Y=15920
X1217 GNDA 13 14 ne3_CDNS_7246548160537 $T=40690 38460 1 0 $X=39890 $Y=27890
X1218 GNDA 13 21 ne3_CDNS_7246548160537 $T=43930 16320 0 0 $X=43130 $Y=15920
X1219 GNDA 13 13 ne3_CDNS_7246548160537 $T=43930 38460 1 0 $X=43130 $Y=27890
X1220 GNDA 13 14 ne3_CDNS_7246548160537 $T=47170 16320 0 0 $X=46370 $Y=15920
X1221 GNDA 13 21 ne3_CDNS_7246548160537 $T=47170 38460 1 0 $X=46370 $Y=27890
X1222 GNDA 13 13 ne3_CDNS_7246548160537 $T=50410 16320 0 0 $X=49610 $Y=15920
X1223 GNDA 13 14 ne3_CDNS_7246548160537 $T=50410 38460 1 0 $X=49610 $Y=27890
X1224 GNDA GNDA GNDA ne3_CDNS_7246548160537 $T=53650 16320 0 0 $X=52850 $Y=15920
X1225 GNDA GNDA GNDA ne3_CDNS_7246548160537 $T=53650 38460 1 0 $X=52850 $Y=27890
X1226 VDDA pe3_CDNS_7246548160538 $T=205435 52315 1 0 $X=203925 $Y=49285
X1227 VDDA pe3_CDNS_7246548160538 $T=205435 175915 1 0 $X=203925 $Y=172885
X1228 VDDA pe3_CDNS_7246548160538 $T=216675 52315 1 0 $X=215165 $Y=49285
X1229 VDDA pe3_CDNS_7246548160538 $T=216675 175915 1 0 $X=215165 $Y=172885
X1230 VDDA pe3_CDNS_7246548160538 $T=227915 52315 1 0 $X=226405 $Y=49285
X1231 VDDA pe3_CDNS_7246548160538 $T=227915 175915 1 0 $X=226405 $Y=172885
X1232 VDDA pe3_CDNS_7246548160538 $T=239155 52315 1 0 $X=237645 $Y=49285
X1233 VDDA pe3_CDNS_7246548160538 $T=239155 175915 1 0 $X=237645 $Y=172885
X1234 VDDA pe3_CDNS_7246548160538 $T=250395 52315 1 0 $X=248885 $Y=49285
X1235 VDDA pe3_CDNS_7246548160538 $T=250395 175915 1 0 $X=248885 $Y=172885
X1236 VDDA pe3_CDNS_7246548160538 $T=261635 52315 1 0 $X=260125 $Y=49285
X1237 VDDA pe3_CDNS_7246548160538 $T=261635 175915 1 0 $X=260125 $Y=172885
X1238 VDDA pe3_CDNS_7246548160538 $T=272875 52315 1 0 $X=271365 $Y=49285
X1239 VDDA pe3_CDNS_7246548160538 $T=272875 175915 1 0 $X=271365 $Y=172885
X1240 VDDA pe3_CDNS_7246548160538 $T=284115 52315 1 0 $X=282605 $Y=49285
X1241 VDDA pe3_CDNS_7246548160538 $T=284115 175915 1 0 $X=282605 $Y=172885
X1242 VDDA pe3_CDNS_7246548160538 $T=295355 52315 1 0 $X=293845 $Y=49285
X1243 VDDA pe3_CDNS_7246548160538 $T=295355 175915 1 0 $X=293845 $Y=172885
X1244 VDDA pe3_CDNS_7246548160538 $T=306595 52315 1 0 $X=305085 $Y=49285
X1245 VDDA pe3_CDNS_7246548160538 $T=306595 175915 1 0 $X=305085 $Y=172885
X1246 VDDA pe3_CDNS_7246548160538 $T=317835 52315 1 0 $X=316325 $Y=49285
X1247 VDDA pe3_CDNS_7246548160538 $T=317835 175915 1 0 $X=316325 $Y=172885
X1248 VDDA pe3_CDNS_7246548160538 $T=329075 52315 1 0 $X=327565 $Y=49285
X1249 VDDA pe3_CDNS_7246548160538 $T=329075 175915 1 0 $X=327565 $Y=172885
X1250 VDDA pe3_CDNS_7246548160538 $T=340315 52315 1 0 $X=338805 $Y=49285
X1251 VDDA pe3_CDNS_7246548160538 $T=340315 175915 1 0 $X=338805 $Y=172885
X1252 VDDA pe3_CDNS_7246548160538 $T=351555 52315 1 0 $X=350045 $Y=49285
X1253 VDDA pe3_CDNS_7246548160538 $T=351555 175915 1 0 $X=350045 $Y=172885
X1254 VDDA pe3_CDNS_7246548160538 $T=362795 52315 1 0 $X=361285 $Y=49285
X1255 VDDA pe3_CDNS_7246548160538 $T=362795 175915 1 0 $X=361285 $Y=172885
X1256 GNDA 25 13 ne3_CDNS_7246548160539 $T=96785 56345 0 0 $X=95985 $Y=55765
X1257 GNDA 25 VOUT ne3_CDNS_7246548160539 $T=102390 56345 0 0 $X=101590 $Y=55765
X1258 VDDA VDDA VDDA 17 16 16 17 MASCO__A15 $T=54830 160530 0 0 $X=54830 $Y=160530
X1259 16 16 VDDA 17 16 16 17 MASCO__A15 $T=99790 160530 0 0 $X=99790 $Y=160530
X1260 VDDA VDDA VDDA 26 17 27 27 MASCO__A15 $T=203925 60085 0 0 $X=203925 $Y=60085
X1261 VDDA VDDA VDDA 26 17 27 28 MASCO__A15 $T=203925 78885 0 0 $X=203925 $Y=78885
X1262 VDDA VDDA VDDA 26 17 27 28 MASCO__A15 $T=203925 97685 0 0 $X=203925 $Y=97685
X1263 VDDA VDDA VDDA 26 17 27 28 MASCO__A15 $T=203925 116485 0 0 $X=203925 $Y=116485
X1264 VDDA VDDA VDDA 26 17 27 28 MASCO__A15 $T=203925 135285 0 0 $X=203925 $Y=135285
X1265 VDDA VDDA VDDA 26 17 26 26 MASCO__A15 $T=203925 154085 0 0 $X=203925 $Y=154085
X1266 27 17 VDDA 27 17 30 26 MASCO__A15 $T=248885 60085 0 0 $X=248885 $Y=60085
X1267 30 17 VDDA 31 17 31 30 MASCO__A15 $T=248885 78885 0 0 $X=248885 $Y=78885
X1268 29 17 VDDA 30 17 24 30 MASCO__A15 $T=248885 97685 0 0 $X=248885 $Y=97685
X1269 30 17 VDDA 29 17 30 28 MASCO__A15 $T=248885 116485 0 0 $X=248885 $Y=116485
X1270 30 17 VDDA 31 17 31 30 MASCO__A15 $T=248885 135285 0 0 $X=248885 $Y=135285
X1271 26 17 VDDA 26 17 27 27 MASCO__A15 $T=248885 154085 0 0 $X=248885 $Y=154085
X1272 26 17 VDDA VDDA VDDA VDDA VDDA MASCO__A15 $T=293845 60085 0 0 $X=293845 $Y=60085
X1273 28 17 VDDA 27 17 26 26 MASCO__A15 $T=293845 78885 0 0 $X=293845 $Y=78885
X1274 28 17 VDDA 27 17 26 26 MASCO__A15 $T=293845 97685 0 0 $X=293845 $Y=97685
X1275 27 17 VDDA 27 17 26 26 MASCO__A15 $T=293845 116485 0 0 $X=293845 $Y=116485
X1276 28 17 VDDA 27 17 26 26 MASCO__A15 $T=293845 135285 0 0 $X=293845 $Y=135285
X1277 27 17 VDDA 30 17 26 26 MASCO__A15 $T=293845 154085 0 0 $X=293845 $Y=154085
D0 GNDA VDDA p_dnw AREA=7.95604e-10 PJ=0.00014876 perimeter=0.00014876 $X=8500 $Y=140710 $dt=6
D1 GNDA VDDA p_dnw AREA=2.14716e-09 PJ=0.0003306 perimeter=0.0003306 $X=48630 $Y=140710 $dt=6
D2 GNDA VDDA p_dnw AREA=3.11448e-11 PJ=3.188e-05 perimeter=3.188e-05 $X=88435 $Y=59745 $dt=6
D3 GNDA 18 p_dnw AREA=1.97548e-10 PJ=8.944e-05 perimeter=8.944e-05 $X=151005 $Y=72505 $dt=6
D4 GNDA 19 p_dnw AREA=1.97548e-10 PJ=8.944e-05 perimeter=8.944e-05 $X=151005 $Y=93985 $dt=6
D5 GNDA 20 p_dnw AREA=1.97548e-10 PJ=8.944e-05 perimeter=8.944e-05 $X=151005 $Y=114935 $dt=6
D6 GNDA VDDA p_dnw AREA=1.47356e-08 PJ=0.0006944 perimeter=0.0006944 $X=181765 $Y=46865 $dt=6
D7 GNDA VDDA p_dnw AREA=1.65707e-09 PJ=0.00035483 perimeter=0.00035483 $X=220785 $Y=22870 $dt=6
D8 GNDA VDDA p_dnw AREA=6.02548e-10 PJ=0.00014223 perimeter=0.00014223 $X=303405 $Y=4665 $dt=6
D9 GNDA VDDA p_ddnw AREA=1.72778e-09 PJ=0.0002104 perimeter=0.0002104 $X=65040 $Y=95265 $dt=7
D10 22 VDDA p_dipdnwmv AREA=9.7703e-10 PJ=0.0001796 perimeter=0.0001796 $X=68890 $Y=99115 $dt=8
D11 GNDA VDDA p_dnw3 AREA=2.92576e-10 PJ=0 perimeter=0 $X=14200 $Y=147550 $dt=9
D12 GNDA VDDA p_dnw3 AREA=2.92576e-10 PJ=0 perimeter=0 $X=14200 $Y=160530 $dt=9
D13 GNDA VDDA p_dnw3 AREA=1.37701e-09 PJ=0 perimeter=0 $X=54830 $Y=147550 $dt=9
D14 GNDA VDDA p_dnw3 AREA=1.37701e-09 PJ=0 perimeter=0 $X=54830 $Y=160530 $dt=9
D15 GNDA VDDA p_dnw3 AREA=2.67592e-11 PJ=0 perimeter=0 $X=89575 $Y=60885 $dt=9
D16 GNDA 18 p_dnw3 AREA=2.77621e-10 PJ=0 perimeter=0 $X=153165 $Y=75665 $dt=9
D17 GNDA 19 p_dnw3 AREA=2.77621e-10 PJ=0 perimeter=0 $X=153165 $Y=97145 $dt=9
D18 GNDA 20 p_dnw3 AREA=2.77621e-10 PJ=0 perimeter=0 $X=153165 $Y=118095 $dt=9
D19 GNDA VDDA p_dnw3 AREA=6.91743e-10 PJ=0 perimeter=0 $X=203925 $Y=49285 $dt=9
D20 GNDA VDDA p_dnw3 AREA=2.05478e-09 PJ=0 perimeter=0 $X=203925 $Y=60085 $dt=9
D21 GNDA VDDA p_dnw3 AREA=2.05478e-09 PJ=0 perimeter=0 $X=203925 $Y=78885 $dt=9
D22 GNDA VDDA p_dnw3 AREA=2.05478e-09 PJ=0 perimeter=0 $X=203925 $Y=97685 $dt=9
D23 GNDA VDDA p_dnw3 AREA=2.05478e-09 PJ=0 perimeter=0 $X=203925 $Y=116485 $dt=9
D24 GNDA VDDA p_dnw3 AREA=2.05478e-09 PJ=0 perimeter=0 $X=203925 $Y=135285 $dt=9
D25 GNDA VDDA p_dnw3 AREA=2.05478e-09 PJ=0 perimeter=0 $X=203925 $Y=154085 $dt=9
D26 GNDA VDDA p_dnw3 AREA=6.91743e-10 PJ=0 perimeter=0 $X=203925 $Y=172885 $dt=9
D27 GNDA VDDA p_dnw3 AREA=2.15633e-10 PJ=0 perimeter=0 $X=222425 $Y=25290 $dt=9
D28 GNDA VDDA p_dnw3 AREA=6.24226e-10 PJ=0 perimeter=0 $X=245245 $Y=25290 $dt=9
D29 GNDA VDDA p_dnw3 AREA=3.27067e-10 PJ=0 perimeter=0 $X=301060 $Y=25290 $dt=9
D30 GNDA VDDA p_dnw3 AREA=5.13756e-11 PJ=0 perimeter=0 $X=305565 $Y=6305 $dt=9
D31 GNDA VDDA p_dnw3 AREA=5.13756e-11 PJ=0 perimeter=0 $X=314825 $Y=6305 $dt=9
D32 GNDA VDDA p_dnw3 AREA=5.13756e-11 PJ=0 perimeter=0 $X=324085 $Y=6305 $dt=9
D33 GNDA VDDA p_dnw3 AREA=1.78488e-10 PJ=0 perimeter=0 $X=331825 $Y=25290 $dt=9
D34 GNDA VDDA p_dnw3 AREA=5.13756e-11 PJ=0 perimeter=0 $X=333345 $Y=6305 $dt=9
D35 GNDA VDDA p_dnw3 AREA=5.13756e-11 PJ=0 perimeter=0 $X=342605 $Y=6305 $dt=9
D36 GNDA VDDA p_dnw3 AREA=1.04198e-10 PJ=0 perimeter=0 $X=350290 $Y=25290 $dt=9
D37 GNDA VDDA p_dnw3 AREA=5.13756e-11 PJ=0 perimeter=0 $X=351865 $Y=6305 $dt=9
D38 GNDA VDDA p_dnw3 AREA=6.70536e-11 PJ=0 perimeter=0 $X=362625 $Y=25290 $dt=9
D39 GNDA VDDA p_dnw3 AREA=4.84812e-11 PJ=0 perimeter=0 $X=372000 $Y=25290 $dt=9
.ends dac6b_amp_n2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pulse_generator                                 *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pulse_generator BIAS1 BIAS2 CUR_OUT D<0> D<1> D<2> D<3> D<4> D<5> ENABLE
+ EXT_FB_RES GNDA GNDHV PULSE_ACTIVE VDD3A VDDHV VREF VSUBHV
** N=19 EP=18 FDC=594
X7 GNDA VDD3A ENABLE BIAS2 PULSE_ACTIVE 1 EXT_FB_RES VSUBHV GNDHV VDDHV
+ CUR_OUT current_source_gm_10_en_r $T=412080 18790 0 0 $X=416015 $Y=22610
X8 GNDA VDD3A mosvc3_CDNS_7246548160521 $T=21090 101820 0 0 $X=20290 $Y=101390
X9 GNDA VDD3A mosvc3_CDNS_7246548160521 $T=21090 154080 1 0 $X=20290 $Y=128460
X10 GNDA VDD3A mosvc3_CDNS_7246548160521 $T=44090 101820 0 0 $X=43290 $Y=101390
X11 GNDA VDD3A mosvc3_CDNS_7246548160521 $T=44090 154080 1 0 $X=43290 $Y=128460
X12 GNDA VDD3A mosvc3_CDNS_7246548160522 $T=422175 183935 0 0 $X=421375 $Y=183505
X13 GNDA VDD3A mosvc3_CDNS_7246548160522 $T=445175 183935 0 0 $X=444375 $Y=183505
X14 GNDA VDD3A mosvc3_CDNS_7246548160522 $T=468175 183935 0 0 $X=467375 $Y=183505
X15 GNDA VDD3A mosvc3_CDNS_7246548160522 $T=491175 183935 0 0 $X=490375 $Y=183505
X16 GNDA VDD3A mosvc3_CDNS_7246548160522 $T=514175 183935 0 0 $X=513375 $Y=183505
X17 GNDA VDD3A mosvc3_CDNS_7246548160522 $T=537175 183935 0 0 $X=536375 $Y=183505
X18 GNDA VDD3A mosvc3_CDNS_7246548160522 $T=560175 183935 0 0 $X=559375 $Y=183505
X19 GNDA VDD3A mosvc3_CDNS_7246548160522 $T=583175 183935 0 0 $X=582375 $Y=183505
X20 GNDA VDD3A BIAS1 ENABLE 1 VREF D<5> D<4> D<3> D<2>
+ D<1> D<0> dac6b_amp_n2 $T=14140 23390 0 0 $X=16780 $Y=24625
R0 GNDA VSUBHV 5 $[s_res] $X=675360 $Y=22605 $dt=5
.ends pulse_generator
