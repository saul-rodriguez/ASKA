* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : constant_gm                                  *
* Netlisted  : Mon Aug 26 08:12:02 2024                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(ne3) nem ndiff(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 1 MP(pe3) pem pdiff(D) p1trm(G) pdiff(S) nwtrm(B)
*.DEVTMPLT 2 NE3I_6() nemi_6 ndiff(D) p1trm(G) ndiff(S) pwitrm(B) dnwtrm(NW) bulk(SB)
*.DEVTMPLT 3 D(p_dnw) p_dnw bulk(POS) nwtrm(NEG)
*.DEVTMPLT 4 D(p_ddnw) p_ddnw bulk(POS) dnwtrm(NEG)
*.DEVTMPLT 5 D(p_dipdnwmv) p_dipwmv pwitrm(POS) dnwtrm(NEG)
*.DEVTMPLT 6 D(p_dnw3) p_dnwm bulk(POS) nwtrm(NEG)
*.DEVTMPLT 7 R(rpp1k1_3) rpp1k1_n p1trm(POS) p1trm(NEG) nwtrm(SUB)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NE3I_6                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NE3I_6 D G S B NW SB
.ends NE3I_6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3i_6_CDNS_724652717070                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3i_6_CDNS_724652717070 1 2 3
** N=3 EP=3 FDC=4
X0 1 3 3 1 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=4.8e-12 ps=1.054e-05 pd=2.096e-05 $X=0 $Y=0 $dt=2
X1 3 3 1 1 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=4.8e-12 ad=2.7e-12 ps=2.096e-05 pd=1.054e-05 $X=3040 $Y=0 $dt=2
D2 1 2 p_ddnw AREA=3.07331e-10 PJ=7.576e-05 perimeter=7.576e-05 $X=-6110 $Y=-4940 $dt=4
D3 1 2 p_dipdnwmv AREA=7.49452e-11 PJ=4.496e-05 perimeter=4.496e-05 $X=-2260 $Y=-1090 $dt=5
.ends ne3i_6_CDNS_724652717070

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724652717071                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724652717071 1 2 3
** N=3 EP=3 FDC=2
M0 2 2 1 1 pe3 L=1e-05 W=2e-06 AD=9.6e-13 AS=9.6e-13 PD=4.96e-06 PS=4.96e-06 $X=0 $Y=0 $dt=1
D1 3 1 p_dnw3 AREA=4.57434e-11 PJ=3.138e-05 perimeter=3.138e-05 $X=-910 $Y=-1440 $dt=6
.ends pe3_CDNS_724652717071

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724652717072                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724652717072 1 2 3 4
** N=4 EP=4 FDC=2
M0 3 2 1 4 ne3 L=2.5e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
M1 1 2 3 4 ne3 L=2.5e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=3040 $Y=0 $dt=0
.ends ne3_CDNS_724652717072

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724652717073                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724652717073 1 2 3 4 5
** N=5 EP=5 FDC=3
M0 3 2 1 4 pe3 L=2.5e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=2.5e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=3040 $Y=0 $dt=1
D2 5 4 p_dnw3 AREA=1.03234e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=6
.ends pe3_CDNS_724652717073

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724652717074                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724652717074 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 3 2 1 4 pe3 L=2.5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
D1 5 4 p_dnw3 AREA=6.65712e-11 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=6
.ends pe3_CDNS_724652717074

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724652717075                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724652717075 1 2 3
*.DEVICECLIMB
** N=4 EP=3 FDC=1
M0 3 2 1 1 pe3 L=2.5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_724652717075

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3i_6_CDNS_724652717076                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3i_6_CDNS_724652717076 1 2 3 4 5
** N=5 EP=5 FDC=10
X0 3 4 5 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=4.8e-12 ps=1.054e-05 pd=2.096e-05 $X=0 $Y=0 $dt=2
X1 5 4 3 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=2.7e-12 ps=1.054e-05 pd=1.054e-05 $X=3040 $Y=0 $dt=2
X2 3 4 5 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=2.7e-12 ps=1.054e-05 pd=1.054e-05 $X=6080 $Y=0 $dt=2
X3 5 4 3 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=2.7e-12 ps=1.054e-05 pd=1.054e-05 $X=9120 $Y=0 $dt=2
X4 3 4 5 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=2.7e-12 ps=1.054e-05 pd=1.054e-05 $X=12160 $Y=0 $dt=2
X5 5 4 3 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=2.7e-12 ps=1.054e-05 pd=1.054e-05 $X=15200 $Y=0 $dt=2
X6 3 4 5 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=2.7e-12 ps=1.054e-05 pd=1.054e-05 $X=18240 $Y=0 $dt=2
X7 5 4 3 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=4.8e-12 ad=2.7e-12 ps=2.096e-05 pd=1.054e-05 $X=21280 $Y=0 $dt=2
D8 1 2 p_ddnw AREA=5.2432e-10 PJ=0.00011224 perimeter=0.00011224 $X=-6110 $Y=-4940 $dt=4
D9 3 2 p_dipdnwmv AREA=1.51486e-10 PJ=8.144e-05 perimeter=8.144e-05 $X=-2260 $Y=-1090 $dt=5
.ends ne3i_6_CDNS_724652717076

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_724652717077                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_724652717077 1 2 3
*.DEVICECLIMB
** N=3 EP=3 FDC=1
R0 2 1 L=0.0002878 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=7
.ends rpp1k1_3_CDNS_724652717077

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: constant_gm                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt constant_gm GNDA OUT1 OUT2 OUT3 VDD3
** N=16 EP=5 FDC=56
X92 GNDA VDD3 5 ne3i_6_CDNS_724652717070 $T=18020 14875 0 0 $X=7250 $Y=5275
X93 15 2 GNDA pe3_CDNS_724652717071 $T=10155 41775 0 0 $X=8645 $Y=39735
X94 4 15 GNDA pe3_CDNS_724652717071 $T=20155 47905 1 180 $X=8645 $Y=45865
X95 5 2 2 GNDA ne3_CDNS_724652717072 $T=25460 39505 0 0 $X=24660 $Y=39105
X96 8 2 4 GNDA ne3_CDNS_724652717072 $T=34790 39505 0 0 $X=33990 $Y=39105
X97 1 4 2 VDD3 GNDA pe3_CDNS_724652717073 $T=11660 58745 0 0 $X=10150 $Y=57715
X98 3 4 4 VDD3 GNDA pe3_CDNS_724652717073 $T=21810 58745 0 0 $X=20300 $Y=57715
X99 7 4 OUT1 VDD3 GNDA pe3_CDNS_724652717073 $T=32565 58745 0 0 $X=31055 $Y=57715
X100 6 4 OUT2 VDD3 GNDA pe3_CDNS_724652717073 $T=43380 58745 0 0 $X=41870 $Y=57715
X101 10 4 OUT3 VDD3 GNDA pe3_CDNS_724652717074 $T=53845 58745 0 0 $X=52335 $Y=57715
X102 VDD3 VDD3 VDD3 pe3_CDNS_724652717075 $T=18765 87600 1 0 $X=17255 $Y=76570
X103 VDD3 VDD3 VDD3 pe3_CDNS_724652717075 $T=18765 106960 1 0 $X=17255 $Y=95930
X104 VDD3 3 6 pe3_CDNS_724652717075 $T=22505 87600 1 0 $X=20995 $Y=76570
X105 VDD3 3 6 pe3_CDNS_724652717075 $T=22505 106960 1 0 $X=20995 $Y=95930
X106 VDD3 3 3 pe3_CDNS_724652717075 $T=26245 87600 1 0 $X=24735 $Y=76570
X107 VDD3 3 1 pe3_CDNS_724652717075 $T=26245 106960 1 0 $X=24735 $Y=95930
X108 VDD3 3 1 pe3_CDNS_724652717075 $T=29985 87600 1 0 $X=28475 $Y=76570
X109 VDD3 3 3 pe3_CDNS_724652717075 $T=29985 106960 1 0 $X=28475 $Y=95930
X110 VDD3 3 7 pe3_CDNS_724652717075 $T=33725 87600 1 0 $X=32215 $Y=76570
X111 VDD3 3 7 pe3_CDNS_724652717075 $T=33725 106960 1 0 $X=32215 $Y=95930
X112 VDD3 VDD3 VDD3 pe3_CDNS_724652717075 $T=37465 87600 1 0 $X=35955 $Y=76570
X113 VDD3 3 10 pe3_CDNS_724652717075 $T=37465 106960 1 0 $X=35955 $Y=95930
X114 VDD3 VDD3 VDD3 pe3_CDNS_724652717075 $T=41205 87600 1 0 $X=39695 $Y=76570
X115 VDD3 VDD3 VDD3 pe3_CDNS_724652717075 $T=41205 106960 1 0 $X=39695 $Y=95930
X116 GNDA VDD3 12 5 8 ne3i_6_CDNS_724652717076 $T=48275 14875 0 0 $X=37505 $Y=5275
X117 GNDA 12 VDD3 rpp1k1_3_CDNS_724652717077 $T=62765 46455 1 90 $X=62545 $Y=41295
D0 GNDA VDD3 p_dnw AREA=4.77568e-10 PJ=0.00014131 perimeter=0.00014131 $X=7700 $Y=53605 $dt=3
D1 GNDA VDD3 p_dnw AREA=1.16854e-09 PJ=0.00017172 perimeter=0.00017172 $X=12555 $Y=74150 $dt=3
D2 GNDA VDD3 p_dnw AREA=1.48411e-09 PJ=0.00019385 perimeter=0.00019385 $X=61625 $Y=40375 $dt=3
D3 GNDA VDD3 p_dnw3 AREA=3.37198e-10 PJ=0 perimeter=0 $X=17255 $Y=76570 $dt=6
D4 GNDA VDD3 p_dnw3 AREA=3.37198e-10 PJ=0 perimeter=0 $X=17255 $Y=95930 $dt=6
.ends constant_gm
