************************************************************************
* auCdl Netlist:
* 
* Library Name:  HVSWITCH
* Top Cell Name: hvswitch5
* View Name:     schematic
* Netlisted on:  Aug  7 16:30:56 2024
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.LDD
*.SCALE METER
.PARAM



************************************************************************
* Library Name: HVSWITCH
* Cell Name:    hvswitch5
* View Name:    schematic
************************************************************************

.SUBCKT hvswitch5 CUR_IN DOWN GNDD GNDHV OUT UP VDD3 VDDHV VSUBHV
*.PININFO CUR_IN:B DOWN:B GNDD:B GNDHV:B OUT:B UP:B VDD3:B VDDHV:B VSUBHV:B
MM4 D4 UPN GNDHV VSUBHV NEDIA W=20u L=1.25u M=1.0 $LDD[NEDIA]
MM2 GATEN DOWNN GNDHV VSUBHV NEDIA W=20u L=1.25u M=1.0 $LDD[NEDIA]
MM0 OUT GATEN CUR_IN VSUBHV NEDIA W=50u L=1.25u M=12.0 $LDD[NEDIA]
RR7 OUT VDDHV 1.00618M $SUB=VSUBHV $[RPP1K1_3] $W=2u $L=2.04358m M=1
RR2 D4 GATEP 125.006K $SUB=VSUBHV $[RPP1K1_3] $W=2u $L=253.7u M=1
RR1 GATEP VDDHV 99.9972K $SUB=VSUBHV $[RPP1K1_3] $W=2u $L=202.9u M=1
RR0 GATEN VDDHV 125.006K $SUB=VSUBHV $[RPP1K1_3] $W=2u $L=253.7u M=1
RR3 GNDHV GATEN 99.9972K $SUB=VSUBHV $[RPP1K1_3] $W=2u $L=202.9u M=1
MM8 UPN net5 GNDD VSUBHV NE3 W=220.0n L=350.0n M=1.0 AD=1.056e-13 AS=1.056e-13 
+ PD=1.4e-06 PS=1.4e-06 NRD=1.22727 NRS=1.22727
MM5 net5 UP GNDD VSUBHV NE3 W=220.0n L=350.0n M=1.0 AD=1.056e-13 AS=1.056e-13 
+ PD=1.4e-06 PS=1.4e-06 NRD=1.22727 NRS=1.22727
MM3 DOWNN DOWN GNDD VSUBHV NE3 W=220.0n L=350.0n M=1.0 AD=1.056e-13 
+ AS=1.056e-13 PD=1.4e-06 PS=1.4e-06 NRD=1.22727 NRS=1.22727
MM7 UPN net5 VDD3 VDD3 PE3 W=440.0n L=300n M=1.0 AD=2.112e-13 AS=2.112e-13 
+ PD=1.84e-06 PS=1.84e-06 NRD=0.613636 NRS=0.613636
MM6 net5 UP VDD3 VDD3 PE3 W=440.0n L=300n M=1.0 AD=2.112e-13 AS=2.112e-13 
+ PD=1.84e-06 PS=1.84e-06 NRD=0.613636 NRS=0.613636
MM11 DOWNN DOWN VDD3 VDD3 PE3 W=440.0n L=300n M=1.0 AD=2.112e-13 AS=2.112e-13 
+ PD=1.84e-06 PS=1.84e-06 NRD=0.613636 NRS=0.613636
MM1 OUT GATEP VDDHV VSUBHV PED W=50u L=940.0n M=12.0 $LDD[PED]
CC2 GNDHV GATEN $[CSF4A] area=6.3936e-11 perimeter=33.72u M=70
CC0 VDDHV OUT $[CSF4A] area=6.3936e-11 perimeter=33.72u M=150
CC4 VDDHV OUT $[CSF4A] area=6.3936e-11 perimeter=33.72u M=150
DD0 GNDHV GATEN DSBA 1.41e-11 3.188e-05 $SUB=VSUBHV M=20.0
DD1 OUT VDDHV DPP20 2.5e-10 110.00000u M=2
.ENDS

