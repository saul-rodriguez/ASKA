* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : ref_bias                                     *
* Netlisted  : Mon Aug 26 08:30:34 2024                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(ne3) nem ndiff(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 1 MP(pe3) pem pdiff(D) p1trm(G) pdiff(S) nwtrm(B)
*.DEVTMPLT 2 NE3I_6() nemi_6 ndiff(D) p1trm(G) ndiff(S) pwitrm(B) dnwtrm(NW) bulk(SB)
*.DEVTMPLT 3 MOSVC3() mosvcm p1trm(G) nwtrm(NW) bulk(SB)
*.DEVTMPLT 4 D(p_dnw) p_dnw bulk(POS) nwtrm(NEG)
*.DEVTMPLT 5 D(p_ddnw) p_ddnw bulk(POS) dnwtrm(NEG)
*.DEVTMPLT 6 D(p_dipdnwmv) p_dipwmv pwitrm(POS) dnwtrm(NEG)
*.DEVTMPLT 7 D(p_dnw3) p_dnwm bulk(POS) nwtrm(NEG)
*.DEVTMPLT 8 R(rpp1k1_3) rpp1k1_s p1trm(POS) p1trm(NEG) bulk(SUB)
*.DEVTMPLT 9 C(cmm5t) cmim capm(POS) m4trm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NE3I_6                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NE3I_6 D G S B NW SB
.ends NE3I_6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MOSVC3                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MOSVC3 G NW SB
.ends MOSVC3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724653828770                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724653828770 1 2 3 4 5
** N=5 EP=5 FDC=11
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=1
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=1
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=1
M4 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=6160 $Y=0 $dt=1
M5 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7700 $Y=0 $dt=1
M6 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=9240 $Y=0 $dt=1
M7 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10780 $Y=0 $dt=1
M8 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12320 $Y=0 $dt=1
M9 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=13860 $Y=0 $dt=1
D10 5 4 p_dnw3 AREA=2.15633e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=7
.ends pe3_CDNS_724653828770

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724653828771                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724653828771 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
.ends ne3_CDNS_724653828771

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724653828772                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724653828772 1 2 3 4 5
** N=5 EP=5 FDC=13
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=1
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=1
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=1
M4 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=6160 $Y=0 $dt=1
M5 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7700 $Y=0 $dt=1
M6 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=9240 $Y=0 $dt=1
M7 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10780 $Y=0 $dt=1
M8 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12320 $Y=0 $dt=1
M9 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=13860 $Y=0 $dt=1
M10 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=15400 $Y=0 $dt=1
M11 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=16940 $Y=0 $dt=1
D12 5 4 p_dnw3 AREA=2.52778e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=7
.ends pe3_CDNS_724653828772

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724653828773                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724653828773 1 2 3 4
** N=4 EP=4 FDC=3
M0 2 2 1 3 pe3 L=2e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 2 3 pe3 L=2e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=2540 $Y=0 $dt=1
D2 4 3 p_dnw3 AREA=9.11736e-11 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=7
.ends pe3_CDNS_724653828773

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_724653828774                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_724653828774 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.0005141 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=8
.ends rpp1k1_3_CDNS_724653828774

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724653828775                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724653828775 1 2 3 4
** N=4 EP=4 FDC=8
M0 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
M1 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=2540 $Y=0 $dt=0
M2 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=5080 $Y=0 $dt=0
M3 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7620 $Y=0 $dt=0
M4 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10160 $Y=0 $dt=0
M5 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12700 $Y=0 $dt=0
M6 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=15240 $Y=0 $dt=0
M7 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=17780 $Y=0 $dt=0
.ends ne3_CDNS_724653828775

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724653828779                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724653828779 1 2 3
*.DEVICECLIMB
** N=4 EP=3 FDC=1
M0 3 2 1 1 pe3 L=2e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_724653828779

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A1 1 2 3 4 5
*.DEVICECLIMB
** N=6 EP=5 FDC=2
X0 1 2 3 pe3_CDNS_724653828779 $T=1510 1030 0 0 $X=0 $Y=0
X1 1 5 4 pe3_CDNS_724653828779 $T=4750 1030 0 0 $X=3240 $Y=0
.ends MASCO__A1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246538287710                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246538287710 1 2 3
*.DEVICECLIMB
** N=4 EP=3 FDC=1
M0 3 2 1 1 pe3 L=1e-05 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_7246538287710

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A2 1 2 3 4 5
*.DEVICECLIMB
** N=6 EP=5 FDC=2
X0 1 4 2 pe3_CDNS_7246538287710 $T=1510 1030 0 0 $X=0 $Y=0
X1 1 5 3 pe3_CDNS_7246538287710 $T=12750 1030 0 0 $X=11240 $Y=0
.ends MASCO__A2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3i_6_CDNS_724653828778                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3i_6_CDNS_724653828778 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=1
X0 1 2 3 1 4 5 NE3I_6 w=1e-05 l=2e-06 as=4.8e-12 ad=4.8e-12 ps=2.096e-05 pd=2.096e-05 $X=0 $Y=0 $dt=2
.ends ne3i_6_CDNS_724653828778

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A3                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A3 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=2
X0 1 4 5 6 7 ne3i_6_CDNS_724653828778 $T=4060 14570 1 0 $X=0 $Y=0
X1 1 2 3 6 7 ne3i_6_CDNS_724653828778 $T=7460 14570 1 0 $X=3400 $Y=0
.ends MASCO__A3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A4                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A4 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=2
X0 1 4 5 6 7 ne3i_6_CDNS_724653828778 $T=4060 4450 0 0 $X=0 $Y=0
X1 1 2 3 6 7 ne3i_6_CDNS_724653828778 $T=7460 4450 0 0 $X=3400 $Y=0
.ends MASCO__A4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__B5                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__B5 1 2 3 4 5 6 7 8 9 10
+ 11
*.DEVICECLIMB
** N=11 EP=11 FDC=4
X0 1 10 6 5 3 2 11 MASCO__A3 $T=0 14680 0 0 $X=0 $Y=14680
X1 1 8 7 9 4 2 11 MASCO__A4 $T=0 0 0 0 $X=0 $Y=0
.ends MASCO__B5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A6                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A6 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=8 EP=7 FDC=4
X0 1 2 3 5 4 MASCO__A1 $T=0 0 0 0 $X=0 $Y=0
X1 1 4 6 7 4 MASCO__A1 $T=6480 0 0 0 $X=6480 $Y=0
.ends MASCO__A6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ref_bias                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ref_bias BIAS GNDA OUT1 OUT2 RES_BIAS VDDA VREF
** N=18 EP=7 FDC=187
X555 11 2 OUT1 VDDA GNDA pe3_CDNS_724653828770 $T=189280 150320 0 0 $X=187770 $Y=149290
X556 12 2 OUT2 VDDA GNDA pe3_CDNS_724653828770 $T=213190 150320 0 0 $X=211680 $Y=149290
X557 GNDA GNDA GNDA ne3_CDNS_724653828771 $T=17980 14080 0 0 $X=17180 $Y=13680
X558 GNDA GNDA GNDA ne3_CDNS_724653828771 $T=17980 30170 0 0 $X=17180 $Y=29770
X559 GNDA 1 3 ne3_CDNS_724653828771 $T=24220 14080 0 0 $X=23420 $Y=13680
X560 GNDA 1 1 ne3_CDNS_724653828771 $T=24220 30170 0 0 $X=23420 $Y=29770
X561 GNDA 1 1 ne3_CDNS_724653828771 $T=30460 14080 0 0 $X=29660 $Y=13680
X562 GNDA 1 3 ne3_CDNS_724653828771 $T=30460 30170 0 0 $X=29660 $Y=29770
X563 GNDA 1 2 ne3_CDNS_724653828771 $T=36700 14080 0 0 $X=35900 $Y=13680
X564 GNDA 1 1 ne3_CDNS_724653828771 $T=36700 30170 0 0 $X=35900 $Y=29770
X565 GNDA 1 1 ne3_CDNS_724653828771 $T=42940 14080 0 0 $X=42140 $Y=13680
X566 GNDA 1 3 ne3_CDNS_724653828771 $T=42940 30170 0 0 $X=42140 $Y=29770
X567 GNDA 1 3 ne3_CDNS_724653828771 $T=49180 14080 0 0 $X=48380 $Y=13680
X568 GNDA GNDA GNDA ne3_CDNS_724653828771 $T=49180 30170 0 0 $X=48380 $Y=29770
X569 GNDA GNDA GNDA ne3_CDNS_724653828771 $T=55420 14080 0 0 $X=54620 $Y=13680
X570 GNDA GNDA GNDA ne3_CDNS_724653828771 $T=55420 30170 0 0 $X=54620 $Y=29770
X571 9 2 RES_BIAS VDDA GNDA pe3_CDNS_724653828772 $T=162340 150320 0 0 $X=160830 $Y=149290
X572 VDDA 8 VDDA GNDA pe3_CDNS_724653828773 $T=138060 190125 0 0 $X=136550 $Y=189095
X573 8 2 VDDA GNDA pe3_CDNS_724653828773 $T=147620 190125 0 0 $X=146110 $Y=189095
X574 RES_BIAS 18 GNDA rpp1k1_3_CDNS_724653828774 $T=87870 117335 0 0 $X=82710 $Y=117115
X575 1 BIAS BIAS GNDA ne3_CDNS_724653828775 $T=17545 54415 0 0 $X=16745 $Y=54015
X576 3 BIAS 6 GNDA ne3_CDNS_724653828775 $T=42480 54195 0 0 $X=41680 $Y=53795
X577 VDDA 16 11 VDDA VDDA MASCO__A1 $T=216005 174905 0 0 $X=216005 $Y=174905
X578 VDDA 16 12 VDDA VDDA MASCO__A1 $T=216005 194925 0 0 $X=216005 $Y=194925
X579 VDDA VDDA 15 VDDA 15 MASCO__A2 $T=10500 171290 0 0 $X=10500 $Y=171290
X580 VDDA VDDA 16 VDDA 15 MASCO__A2 $T=10500 188970 0 0 $X=10500 $Y=188970
X581 VDDA 16 15 15 15 MASCO__A2 $T=32980 171290 0 0 $X=32980 $Y=171290
X582 VDDA 15 16 15 15 MASCO__A2 $T=32980 188970 0 0 $X=32980 $Y=188970
X583 VDDA 16 15 15 15 MASCO__A2 $T=55460 171290 0 0 $X=55460 $Y=171290
X584 VDDA 15 16 15 15 MASCO__A2 $T=55460 188970 0 0 $X=55460 $Y=188970
X585 VDDA 16 15 15 15 MASCO__A2 $T=77940 171290 0 0 $X=77940 $Y=171290
X586 VDDA 15 16 15 15 MASCO__A2 $T=77940 188970 0 0 $X=77940 $Y=188970
X587 VDDA 16 VDDA 15 VDDA MASCO__A2 $T=100420 171290 0 0 $X=100420 $Y=171290
X588 VDDA 15 VDDA 15 VDDA MASCO__A2 $T=100420 188970 0 0 $X=100420 $Y=188970
X589 6 VDDA 6 6 6 16 15 RES_BIAS 6 VREF
+ GNDA MASCO__B5 $T=9330 114030 0 0 $X=9330 $Y=114030
X590 6 VDDA 15 16 RES_BIAS 16 15 RES_BIAS VREF VREF
+ GNDA MASCO__B5 $T=16130 114030 0 0 $X=16130 $Y=114030
X591 6 VDDA 15 16 RES_BIAS 16 15 RES_BIAS VREF VREF
+ GNDA MASCO__B5 $T=22930 114030 0 0 $X=22930 $Y=114030
X592 6 VDDA 15 16 RES_BIAS 16 15 RES_BIAS VREF VREF
+ GNDA MASCO__B5 $T=29730 114030 0 0 $X=29730 $Y=114030
X593 6 VDDA 15 16 RES_BIAS 16 15 RES_BIAS VREF VREF
+ GNDA MASCO__B5 $T=36530 114030 0 0 $X=36530 $Y=114030
X594 6 VDDA 15 16 RES_BIAS 16 15 RES_BIAS VREF VREF
+ GNDA MASCO__B5 $T=43330 114030 0 0 $X=43330 $Y=114030
X595 6 VDDA 15 16 RES_BIAS 16 15 RES_BIAS VREF VREF
+ GNDA MASCO__B5 $T=50130 114030 0 0 $X=50130 $Y=114030
X596 6 VDDA 15 16 RES_BIAS 6 6 6 VREF 6
+ GNDA MASCO__B5 $T=56930 114030 0 0 $X=56930 $Y=114030
X597 VDDA VDDA VDDA 16 11 12 9 MASCO__A6 $T=164165 174905 0 0 $X=164165 $Y=174905
X598 VDDA VDDA VDDA 16 12 9 11 MASCO__A6 $T=164165 194925 0 0 $X=164165 $Y=194925
X599 VDDA 16 11 16 9 12 9 MASCO__A6 $T=177125 174905 0 0 $X=177125 $Y=174905
X600 VDDA 16 12 16 12 9 11 MASCO__A6 $T=177125 194925 0 0 $X=177125 $Y=194925
X601 VDDA 16 11 16 9 12 9 MASCO__A6 $T=190085 174905 0 0 $X=190085 $Y=174905
X602 VDDA 16 9 16 12 9 11 MASCO__A6 $T=190085 194925 0 0 $X=190085 $Y=194925
X603 VDDA 16 11 16 11 12 9 MASCO__A6 $T=203045 174905 0 0 $X=203045 $Y=174905
X604 VDDA 16 9 16 12 9 11 MASCO__A6 $T=203045 194925 0 0 $X=203045 $Y=194925
X605 OUT2 GNDA GNDA MOSVC3 w=3e-05 l=3e-05 $X=85530 $Y=8110 $dt=3
X606 OUT2 GNDA GNDA MOSVC3 w=3e-05 l=3e-05 $X=85530 $Y=39350 $dt=3
X607 OUT2 GNDA GNDA MOSVC3 w=3e-05 l=3e-05 $X=85530 $Y=70590 $dt=3
X608 OUT1 GNDA GNDA MOSVC3 w=3e-05 l=3e-05 $X=122495 $Y=8050 $dt=3
X609 OUT1 GNDA GNDA MOSVC3 w=3e-05 l=3e-05 $X=122495 $Y=39290 $dt=3
X610 OUT1 GNDA GNDA MOSVC3 w=3e-05 l=3e-05 $X=122495 $Y=70530 $dt=3
D6 GNDA VDDA p_dnw AREA=2.36318e-09 PJ=0.00033402 perimeter=0.00033402 $X=4385 $Y=163650 $dt=4
D7 GNDA VDDA p_dnw AREA=2.57209e-10 PJ=8.388e-05 perimeter=8.388e-05 $X=134410 $Y=183535 $dt=4
D8 GNDA VDDA p_dnw AREA=1.81014e-09 PJ=0.00023539 perimeter=0.00023539 $X=158410 $Y=166295 $dt=4
D9 GNDA VDDA p_dnw AREA=8.15582e-10 PJ=0.0001871 perimeter=0.0001871 $X=158690 $Y=143730 $dt=4
D10 GNDA VDDA p_dnw AREA=9.45702e-09 PJ=0.00040696 perimeter=0.00040696 $X=159475 $Y=6005 $dt=4
D11 GNDA VDDA p_ddnw AREA=1.66704e-09 PJ=0.0001998 perimeter=0.0001998 $X=8060 $Y=112760 $dt=5
D12 6 VDDA p_dipdnwmv AREA=9.57098e-10 PJ=0.000169 perimeter=0.000169 $X=11910 $Y=116610 $dt=6
D13 GNDA VDDA p_dnw3 AREA=1.37701e-09 PJ=0 perimeter=0 $X=10500 $Y=171290 $dt=7
D14 GNDA VDDA p_dnw3 AREA=1.37701e-09 PJ=0 perimeter=0 $X=10500 $Y=188970 $dt=7
D15 GNDA GNDA p_dnw3 AREA=2.03309e-10 PJ=0.00024988 perimeter=0.00024988 $X=85100 $Y=7310 $dt=7
D16 GNDA GNDA p_dnw3 AREA=2.03309e-10 PJ=0.00024988 perimeter=0.00024988 $X=122065 $Y=7250 $dt=7
D17 GNDA VDDA p_dnw3 AREA=7.24806e-10 PJ=0 perimeter=0 $X=164165 $Y=174905 $dt=7
D18 GNDA VDDA p_dnw3 AREA=7.24806e-10 PJ=0 perimeter=0 $X=164165 $Y=194925 $dt=7
C19 16 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=161615 $Y=8145 $dt=9
C20 16 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=161615 $Y=39745 $dt=9
C21 16 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=161615 $Y=71345 $dt=9
C22 16 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=161615 $Y=102945 $dt=9
C23 16 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=196615 $Y=8145 $dt=9
C24 16 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=196615 $Y=39745 $dt=9
C25 16 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=196615 $Y=71345 $dt=9
C26 16 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=196615 $Y=102945 $dt=9
.ends ref_bias
