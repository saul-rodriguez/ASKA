* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : por2                                         *
* Netlisted  : Mon Aug 26 08:07:33 2024                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(ne3) nem ndiff(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 1 MP(pe3) pem pdiff(D) p1trm(G) pdiff(S) nwtrm(B)
*.DEVTMPLT 2 MOSVC3() mosvcm p1trm(G) nwtrm(NW) bulk(SB)
*.DEVTMPLT 3 D(p_dnw) p_dnw bulk(POS) nwtrm(NEG)
*.DEVTMPLT 4 D(p_dnw3) p_dnwm bulk(POS) nwtrm(NEG)
*.DEVTMPLT 5 R(rpp1k1_3) rpp1k1_s p1trm(POS) p1trm(NEG) bulk(SUB)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_724652447320                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_724652447320 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_724652447320

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_724652447321                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_724652447321 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_724652447321

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_724652447322                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_724652447322 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_724652447322

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724652447323                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724652447323 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724652447323

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724652447324                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724652447324 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724652447324

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724652447325                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724652447325 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724652447325

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724652447326                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724652447326 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724652447326

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_724652447327                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_724652447327 1 2
** N=2 EP=2 FDC=0
.ends VIA2_C_CDNS_724652447327

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246524473210                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246524473210 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246524473210

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: STE_3VX4                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt STE_3VX4 1 2 3 4
** N=7 EP=4 FDC=15
M0 5 3 6 2 ne3 L=3.5e-07 W=7.6e-07 AD=2.15279e-13 AS=3.648e-13 PD=1.40142e-06 PS=2.48e-06 $X=620 $Y=660 $dt=0
M1 2 3 5 2 ne3 L=3.5e-07 W=6.5e-07 AD=5.1e-13 AS=1.84121e-13 PD=3.09e-06 PS=1.19858e-06 $X=1510 $Y=660 $dt=0
M2 1 6 5 2 ne3 L=3.5e-07 W=8.9e-07 AD=4.628e-13 AS=5.162e-13 PD=2.82e-06 PS=2.94e-06 $X=3790 $Y=660 $dt=0
M3 4 6 2 2 ne3 L=3.5e-07 W=6.6e-07 AD=1.782e-13 AS=5.8405e-13 PD=1.2e-06 PS=3.57e-06 $X=6040 $Y=865 $dt=0
M4 2 6 4 2 ne3 L=3.5e-07 W=6.6e-07 AD=3.2115e-13 AS=1.782e-13 PD=1.835e-06 PS=1.2e-06 $X=6930 $Y=865 $dt=0
M5 4 6 2 2 ne3 L=3.5e-07 W=6.6e-07 AD=1.782e-13 AS=3.2115e-13 PD=1.2e-06 PS=1.835e-06 $X=7900 $Y=865 $dt=0
M6 2 6 4 2 ne3 L=3.5e-07 W=6.6e-07 AD=6.249e-13 AS=1.782e-13 PD=3.55e-06 PS=1.2e-06 $X=8790 $Y=865 $dt=0
M7 7 3 6 1 pe3 L=3e-07 W=1.41e-06 AD=4.21161e-13 AS=7.1205e-13 PD=2.04348e-06 PS=3.83e-06 $X=645 $Y=2410 $dt=1
M8 1 3 7 1 pe3 L=3e-07 W=1.35e-06 AD=9.5195e-13 AS=4.03239e-13 PD=4.66e-06 PS=1.95652e-06 $X=1535 $Y=2410 $dt=1
M9 2 6 7 1 pe3 L=3.5e-07 W=1.41e-06 AD=6.768e-13 AS=8.178e-13 PD=3.78e-06 PS=3.98e-06 $X=3790 $Y=2410 $dt=1
M10 4 6 1 1 pe3 L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=9.5945e-13 PD=2e-06 PS=4.66e-06 $X=6145 $Y=2410 $dt=1
M11 1 6 4 1 pe3 L=3e-07 W=1.41e-06 AD=4.1765e-13 AS=4.1595e-13 PD=2.01e-06 PS=2e-06 $X=7035 $Y=2410 $dt=1
M12 4 6 1 1 pe3 L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=4.1765e-13 PD=2e-06 PS=2.01e-06 $X=7925 $Y=2410 $dt=1
M13 1 6 4 1 pe3 L=3e-07 W=1.41e-06 AD=9.8585e-13 AS=4.1595e-13 PD=4.69e-06 PS=2e-06 $X=8815 $Y=2410 $dt=1
D14 2 1 p_dnw3 AREA=3.43516e-11 PJ=2.816e-05 perimeter=2.816e-05 $X=-430 $Y=1980 $dt=4
.ends STE_3VX4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724652447320                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724652447320 1 2 3
** N=3 EP=3 FDC=2
M0 3 2 1 1 ne3 L=3.5e-07 W=5e-06 AD=1.35e-12 AS=2.4e-12 PD=5.54e-06 PS=1.096e-05 $X=0 $Y=0 $dt=0
M1 1 2 3 1 ne3 L=3.5e-07 W=5e-06 AD=2.4e-12 AS=1.35e-12 PD=1.096e-05 PS=5.54e-06 $X=890 $Y=0 $dt=0
.ends ne3_CDNS_724652447320

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724652447322                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724652447322 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=5e-06 W=5e-06 AD=2.4e-12 AS=2.4e-12 PD=1.096e-05 PS=1.096e-05 $X=0 $Y=0 $dt=0
.ends ne3_CDNS_724652447322

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724652447323                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724652447323 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=1
M0 3 2 1 4 pe3 L=5e-07 W=4e-06 AD=1.92e-12 AS=1.92e-12 PD=8.96e-06 PS=8.96e-06 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_724652447323

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_724652447324                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_724652447324 1 2
** N=2 EP=2 FDC=1
R0 2 1 L=0.00283888 W=4e-06 $[rpp1k1_3] $SUB=1 $X=-4220 $Y=0 $dt=5
.ends rpp1k1_3_CDNS_724652447324

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_724652447327                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_724652447327 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.00411438 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=5
.ends rpp1k1_3_CDNS_724652447327

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724652447326                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724652447326 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
M0 3 2 1 1 pe3 L=5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_724652447326

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A1 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 2 3 6 pe3_CDNS_724652447326 $T=1510 1030 0 0 $X=0 $Y=0
X1 1 4 5 6 pe3_CDNS_724652447326 $T=7750 1030 0 0 $X=6240 $Y=0
.ends MASCO__A1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724652447321                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724652447321 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
.ends ne3_CDNS_724652447321

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A2 1 2 3 4
** N=4 EP=4 FDC=2
X0 1 2 2 ne3_CDNS_724652447321 $T=800 400 0 0 $X=0 $Y=0
X1 1 4 3 ne3_CDNS_724652447321 $T=7040 400 0 0 $X=6240 $Y=0
.ends MASCO__A2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: por2                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt por2 9 1 2 11 3
** N=11 EP=5 FDC=95
X0 1 VIA2_C_CDNS_724652447320 $T=15255 137415 0 0 $X=14285 $Y=136755
X1 1 VIA2_C_CDNS_724652447320 $T=15255 152405 0 0 $X=14285 $Y=151745
X2 1 VIA2_C_CDNS_724652447320 $T=15255 167375 0 0 $X=14285 $Y=166715
X3 2 VIA2_C_CDNS_724652447320 $T=17595 139255 0 0 $X=16625 $Y=138595
X4 2 VIA2_C_CDNS_724652447320 $T=17595 154245 0 0 $X=16625 $Y=153585
X5 2 VIA2_C_CDNS_724652447320 $T=70555 139255 0 0 $X=69585 $Y=138595
X6 2 VIA2_C_CDNS_724652447320 $T=70555 154245 0 0 $X=69585 $Y=153585
X7 1 VIA2_C_CDNS_724652447320 $T=72895 137415 0 0 $X=71925 $Y=136755
X8 1 VIA2_C_CDNS_724652447320 $T=72895 152405 0 0 $X=71925 $Y=151745
X9 1 VIA2_C_CDNS_724652447320 $T=72895 167375 0 0 $X=71925 $Y=166715
X10 3 VIA2_C_CDNS_724652447321 $T=23865 178015 0 0 $X=22375 $Y=177615
X11 3 VIA2_C_CDNS_724652447321 $T=23865 195635 0 0 $X=22375 $Y=195235
X12 3 VIA2_C_CDNS_724652447321 $T=23865 213695 0 0 $X=22375 $Y=213295
X13 3 VIA2_C_CDNS_724652447321 $T=23865 231315 0 0 $X=22375 $Y=230915
X14 3 VIA2_C_CDNS_724652447321 $T=91605 178015 0 0 $X=90115 $Y=177615
X15 3 VIA2_C_CDNS_724652447321 $T=91605 195635 0 0 $X=90115 $Y=195235
X16 3 VIA2_C_CDNS_724652447321 $T=91605 213695 0 0 $X=90115 $Y=213295
X17 3 VIA2_C_CDNS_724652447321 $T=91605 231315 0 0 $X=90115 $Y=230915
X18 4 VIA2_C_CDNS_724652447322 $T=19555 176735 0 0 $X=18895 $Y=176285
X19 4 VIA2_C_CDNS_724652447322 $T=19555 194355 0 0 $X=18895 $Y=193905
X20 4 VIA2_C_CDNS_724652447322 $T=19555 212415 0 0 $X=18895 $Y=211965
X21 4 VIA2_C_CDNS_724652447322 $T=19555 230035 0 0 $X=18895 $Y=229585
X22 5 VIA2_C_CDNS_724652447322 $T=21335 175455 0 0 $X=20675 $Y=175005
X23 5 VIA2_C_CDNS_724652447322 $T=21335 193075 0 0 $X=20675 $Y=192625
X24 5 VIA2_C_CDNS_724652447322 $T=21335 211135 0 0 $X=20675 $Y=210685
X25 5 VIA2_C_CDNS_724652447322 $T=21335 228755 0 0 $X=20675 $Y=228305
X26 4 VIA2_C_CDNS_724652447322 $T=94135 176735 0 0 $X=93475 $Y=176285
X27 4 VIA2_C_CDNS_724652447322 $T=94135 194355 0 0 $X=93475 $Y=193905
X28 4 VIA2_C_CDNS_724652447322 $T=94135 212415 0 0 $X=93475 $Y=211965
X29 4 VIA2_C_CDNS_724652447322 $T=94135 230035 0 0 $X=93475 $Y=229585
X30 5 VIA2_C_CDNS_724652447322 $T=95915 175455 0 0 $X=95255 $Y=175005
X31 5 VIA2_C_CDNS_724652447322 $T=95915 193075 0 0 $X=95255 $Y=192625
X32 5 VIA2_C_CDNS_724652447322 $T=95915 211135 0 0 $X=95255 $Y=210685
X33 5 VIA2_C_CDNS_724652447322 $T=95915 228755 0 0 $X=95255 $Y=228305
X34 6 VIA2_C_CDNS_724652447322 $T=97695 191795 0 0 $X=97035 $Y=191345
X35 6 VIA2_C_CDNS_724652447322 $T=97695 209855 0 0 $X=97035 $Y=209405
X36 6 VIA2_C_CDNS_724652447322 $T=97695 227475 0 0 $X=97035 $Y=227025
X37 3 VIA1_C_CDNS_724652447323 $T=26885 178015 0 0 $X=26745 $Y=177565
X38 3 VIA1_C_CDNS_724652447323 $T=26885 195635 0 0 $X=26745 $Y=195185
X39 3 VIA1_C_CDNS_724652447323 $T=26885 213695 0 0 $X=26745 $Y=213245
X40 3 VIA1_C_CDNS_724652447323 $T=29655 195635 0 0 $X=29515 $Y=195185
X41 3 VIA1_C_CDNS_724652447323 $T=29655 213695 0 0 $X=29515 $Y=213245
X42 3 VIA1_C_CDNS_724652447323 $T=29655 231315 0 0 $X=29515 $Y=230865
X43 3 VIA1_C_CDNS_724652447323 $T=32425 178015 0 0 $X=32285 $Y=177565
X44 3 VIA1_C_CDNS_724652447323 $T=32425 195635 0 0 $X=32285 $Y=195185
X45 3 VIA1_C_CDNS_724652447323 $T=32425 213695 0 0 $X=32285 $Y=213245
X46 3 VIA1_C_CDNS_724652447323 $T=33125 178015 0 0 $X=32985 $Y=177565
X47 3 VIA1_C_CDNS_724652447323 $T=33125 195635 0 0 $X=32985 $Y=195185
X48 3 VIA1_C_CDNS_724652447323 $T=33125 213695 0 0 $X=32985 $Y=213245
X49 5 VIA1_C_CDNS_724652447323 $T=35895 193075 0 0 $X=35755 $Y=192625
X50 5 VIA1_C_CDNS_724652447323 $T=35895 211135 0 0 $X=35755 $Y=210685
X51 5 VIA1_C_CDNS_724652447323 $T=35895 228755 0 0 $X=35755 $Y=228305
X52 4 VIA1_C_CDNS_724652447323 $T=38665 176735 0 0 $X=38525 $Y=176285
X53 5 VIA1_C_CDNS_724652447323 $T=38665 193075 0 0 $X=38525 $Y=192625
X54 4 VIA1_C_CDNS_724652447323 $T=38665 212415 0 0 $X=38525 $Y=211965
X55 3 VIA1_C_CDNS_724652447323 $T=39365 178015 0 0 $X=39225 $Y=177565
X56 3 VIA1_C_CDNS_724652447323 $T=39365 195635 0 0 $X=39225 $Y=195185
X57 3 VIA1_C_CDNS_724652447323 $T=39365 213695 0 0 $X=39225 $Y=213245
X58 5 VIA1_C_CDNS_724652447323 $T=42135 193075 0 0 $X=41995 $Y=192625
X59 5 VIA1_C_CDNS_724652447323 $T=42135 211135 0 0 $X=41995 $Y=210685
X60 5 VIA1_C_CDNS_724652447323 $T=42135 228755 0 0 $X=41995 $Y=228305
X61 5 VIA1_C_CDNS_724652447323 $T=44905 175455 0 0 $X=44765 $Y=175005
X62 4 VIA1_C_CDNS_724652447323 $T=44905 194355 0 0 $X=44765 $Y=193905
X63 5 VIA1_C_CDNS_724652447323 $T=44905 211135 0 0 $X=44765 $Y=210685
X64 3 VIA1_C_CDNS_724652447323 $T=45605 178015 0 0 $X=45465 $Y=177565
X65 3 VIA1_C_CDNS_724652447323 $T=45605 195635 0 0 $X=45465 $Y=195185
X66 3 VIA1_C_CDNS_724652447323 $T=45605 213695 0 0 $X=45465 $Y=213245
X67 5 VIA1_C_CDNS_724652447323 $T=48375 193075 0 0 $X=48235 $Y=192625
X68 5 VIA1_C_CDNS_724652447323 $T=48375 211135 0 0 $X=48235 $Y=210685
X69 5 VIA1_C_CDNS_724652447323 $T=48375 228755 0 0 $X=48235 $Y=228305
X70 4 VIA1_C_CDNS_724652447323 $T=51145 176735 0 0 $X=51005 $Y=176285
X71 6 VIA1_C_CDNS_724652447323 $T=51145 191795 0 0 $X=51005 $Y=191345
X72 4 VIA1_C_CDNS_724652447323 $T=51145 212415 0 0 $X=51005 $Y=211965
X73 3 VIA1_C_CDNS_724652447323 $T=51845 178015 0 0 $X=51705 $Y=177565
X74 3 VIA1_C_CDNS_724652447323 $T=51845 195635 0 0 $X=51705 $Y=195185
X75 3 VIA1_C_CDNS_724652447323 $T=51845 213695 0 0 $X=51705 $Y=213245
X76 5 VIA1_C_CDNS_724652447323 $T=54615 193075 0 0 $X=54475 $Y=192625
X77 5 VIA1_C_CDNS_724652447323 $T=54615 211135 0 0 $X=54475 $Y=210685
X78 5 VIA1_C_CDNS_724652447323 $T=54615 228755 0 0 $X=54475 $Y=228305
X79 5 VIA1_C_CDNS_724652447323 $T=57385 175455 0 0 $X=57245 $Y=175005
X80 4 VIA1_C_CDNS_724652447323 $T=57385 194355 0 0 $X=57245 $Y=193905
X81 5 VIA1_C_CDNS_724652447323 $T=57385 211135 0 0 $X=57245 $Y=210685
X82 3 VIA1_C_CDNS_724652447323 $T=58085 178015 0 0 $X=57945 $Y=177565
X83 3 VIA1_C_CDNS_724652447323 $T=58085 195635 0 0 $X=57945 $Y=195185
X84 3 VIA1_C_CDNS_724652447323 $T=58085 213695 0 0 $X=57945 $Y=213245
X85 5 VIA1_C_CDNS_724652447323 $T=60855 193075 0 0 $X=60715 $Y=192625
X86 5 VIA1_C_CDNS_724652447323 $T=60855 211135 0 0 $X=60715 $Y=210685
X87 5 VIA1_C_CDNS_724652447323 $T=60855 228755 0 0 $X=60715 $Y=228305
X88 4 VIA1_C_CDNS_724652447323 $T=63625 176735 0 0 $X=63485 $Y=176285
X89 5 VIA1_C_CDNS_724652447323 $T=63625 193075 0 0 $X=63485 $Y=192625
X90 4 VIA1_C_CDNS_724652447323 $T=63625 212415 0 0 $X=63485 $Y=211965
X91 3 VIA1_C_CDNS_724652447323 $T=64325 178015 0 0 $X=64185 $Y=177565
X92 3 VIA1_C_CDNS_724652447323 $T=64325 195635 0 0 $X=64185 $Y=195185
X93 3 VIA1_C_CDNS_724652447323 $T=64325 213695 0 0 $X=64185 $Y=213245
X94 5 VIA1_C_CDNS_724652447323 $T=67095 193075 0 0 $X=66955 $Y=192625
X95 5 VIA1_C_CDNS_724652447323 $T=67095 211135 0 0 $X=66955 $Y=210685
X96 5 VIA1_C_CDNS_724652447323 $T=67095 228755 0 0 $X=66955 $Y=228305
X97 5 VIA1_C_CDNS_724652447323 $T=69865 175455 0 0 $X=69725 $Y=175005
X98 6 VIA1_C_CDNS_724652447323 $T=69865 191795 0 0 $X=69725 $Y=191345
X99 5 VIA1_C_CDNS_724652447323 $T=69865 211135 0 0 $X=69725 $Y=210685
X100 3 VIA1_C_CDNS_724652447323 $T=70565 178015 0 0 $X=70425 $Y=177565
X101 3 VIA1_C_CDNS_724652447323 $T=70565 195635 0 0 $X=70425 $Y=195185
X102 3 VIA1_C_CDNS_724652447323 $T=70565 213695 0 0 $X=70425 $Y=213245
X103 5 VIA1_C_CDNS_724652447323 $T=73335 193075 0 0 $X=73195 $Y=192625
X104 5 VIA1_C_CDNS_724652447323 $T=73335 211135 0 0 $X=73195 $Y=210685
X105 5 VIA1_C_CDNS_724652447323 $T=73335 228755 0 0 $X=73195 $Y=228305
X106 4 VIA1_C_CDNS_724652447323 $T=76105 176735 0 0 $X=75965 $Y=176285
X107 5 VIA1_C_CDNS_724652447323 $T=76105 193075 0 0 $X=75965 $Y=192625
X108 4 VIA1_C_CDNS_724652447323 $T=76105 212415 0 0 $X=75965 $Y=211965
X109 3 VIA1_C_CDNS_724652447323 $T=76805 178015 0 0 $X=76665 $Y=177565
X110 3 VIA1_C_CDNS_724652447323 $T=76805 195635 0 0 $X=76665 $Y=195185
X111 3 VIA1_C_CDNS_724652447323 $T=76805 213695 0 0 $X=76665 $Y=213245
X112 5 VIA1_C_CDNS_724652447323 $T=79575 193075 0 0 $X=79435 $Y=192625
X113 3 VIA1_C_CDNS_724652447323 $T=79575 213695 0 0 $X=79435 $Y=213245
X114 3 VIA1_C_CDNS_724652447323 $T=79575 231315 0 0 $X=79435 $Y=230865
X115 5 VIA1_C_CDNS_724652447323 $T=82345 175455 0 0 $X=82205 $Y=175005
X116 3 VIA1_C_CDNS_724652447323 $T=82345 195635 0 0 $X=82205 $Y=195185
X117 3 VIA1_C_CDNS_724652447323 $T=82345 213695 0 0 $X=82205 $Y=213245
X118 3 VIA1_C_CDNS_724652447323 $T=83045 178015 0 0 $X=82905 $Y=177565
X119 3 VIA1_C_CDNS_724652447323 $T=83045 195635 0 0 $X=82905 $Y=195185
X120 3 VIA1_C_CDNS_724652447323 $T=83045 213695 0 0 $X=82905 $Y=213245
X121 3 VIA1_C_CDNS_724652447323 $T=85815 195635 0 0 $X=85675 $Y=195185
X122 3 VIA1_C_CDNS_724652447323 $T=85815 213695 0 0 $X=85675 $Y=213245
X123 3 VIA1_C_CDNS_724652447323 $T=85815 231315 0 0 $X=85675 $Y=230865
X124 3 VIA1_C_CDNS_724652447323 $T=88585 178015 0 0 $X=88445 $Y=177565
X125 3 VIA1_C_CDNS_724652447323 $T=88585 195635 0 0 $X=88445 $Y=195185
X126 3 VIA1_C_CDNS_724652447323 $T=88585 213695 0 0 $X=88445 $Y=213245
X127 2 VIA1_C_CDNS_724652447324 $T=19465 139255 0 0 $X=19325 $Y=138545
X128 2 VIA1_C_CDNS_724652447324 $T=19465 154245 0 0 $X=19325 $Y=153535
X129 2 VIA1_C_CDNS_724652447324 $T=25005 139255 0 0 $X=24865 $Y=138545
X130 2 VIA1_C_CDNS_724652447324 $T=25005 154245 0 0 $X=24865 $Y=153535
X131 2 VIA1_C_CDNS_724652447324 $T=25705 139255 0 0 $X=25565 $Y=138545
X132 2 VIA1_C_CDNS_724652447324 $T=25705 154245 0 0 $X=25565 $Y=153535
X133 1 VIA1_C_CDNS_724652447324 $T=28475 152405 0 0 $X=28335 $Y=151695
X134 1 VIA1_C_CDNS_724652447324 $T=28475 167375 0 0 $X=28335 $Y=166665
X135 1 VIA1_C_CDNS_724652447324 $T=31245 137415 0 0 $X=31105 $Y=136705
X136 1 VIA1_C_CDNS_724652447324 $T=31245 152405 0 0 $X=31105 $Y=151695
X137 2 VIA1_C_CDNS_724652447324 $T=31945 139255 0 0 $X=31805 $Y=138545
X138 2 VIA1_C_CDNS_724652447324 $T=31945 154245 0 0 $X=31805 $Y=153535
X139 1 VIA1_C_CDNS_724652447324 $T=34715 152405 0 0 $X=34575 $Y=151695
X140 1 VIA1_C_CDNS_724652447324 $T=34715 167375 0 0 $X=34575 $Y=166665
X141 1 VIA1_C_CDNS_724652447324 $T=37485 137415 0 0 $X=37345 $Y=136705
X142 1 VIA1_C_CDNS_724652447324 $T=37485 152405 0 0 $X=37345 $Y=151695
X143 2 VIA1_C_CDNS_724652447324 $T=38185 139255 0 0 $X=38045 $Y=138545
X144 2 VIA1_C_CDNS_724652447324 $T=38185 154245 0 0 $X=38045 $Y=153535
X145 1 VIA1_C_CDNS_724652447324 $T=40955 152405 0 0 $X=40815 $Y=151695
X146 1 VIA1_C_CDNS_724652447324 $T=40955 167375 0 0 $X=40815 $Y=166665
X147 5 VIA1_C_CDNS_724652447324 $T=43725 135575 0 0 $X=43585 $Y=134865
X148 1 VIA1_C_CDNS_724652447324 $T=43725 152405 0 0 $X=43585 $Y=151695
X149 2 VIA1_C_CDNS_724652447324 $T=44425 139255 0 0 $X=44285 $Y=138545
X150 2 VIA1_C_CDNS_724652447324 $T=44425 154245 0 0 $X=44285 $Y=153535
X151 1 VIA1_C_CDNS_724652447324 $T=47195 152405 0 0 $X=47055 $Y=151695
X152 1 VIA1_C_CDNS_724652447324 $T=47195 167375 0 0 $X=47055 $Y=166665
X153 1 VIA1_C_CDNS_724652447324 $T=49965 137415 0 0 $X=49825 $Y=136705
X154 1 VIA1_C_CDNS_724652447324 $T=49965 152405 0 0 $X=49825 $Y=151695
X155 2 VIA1_C_CDNS_724652447324 $T=50665 139255 0 0 $X=50525 $Y=138545
X156 2 VIA1_C_CDNS_724652447324 $T=50665 154245 0 0 $X=50525 $Y=153535
X157 1 VIA1_C_CDNS_724652447324 $T=53435 152405 0 0 $X=53295 $Y=151695
X158 1 VIA1_C_CDNS_724652447324 $T=53435 167375 0 0 $X=53295 $Y=166665
X159 1 VIA1_C_CDNS_724652447324 $T=56205 137415 0 0 $X=56065 $Y=136705
X160 1 VIA1_C_CDNS_724652447324 $T=56205 152405 0 0 $X=56065 $Y=151695
X161 2 VIA1_C_CDNS_724652447324 $T=56905 139255 0 0 $X=56765 $Y=138545
X162 2 VIA1_C_CDNS_724652447324 $T=56905 154245 0 0 $X=56765 $Y=153535
X163 1 VIA1_C_CDNS_724652447324 $T=59675 152405 0 0 $X=59535 $Y=151695
X164 1 VIA1_C_CDNS_724652447324 $T=62445 137415 0 0 $X=62305 $Y=136705
X165 2 VIA1_C_CDNS_724652447324 $T=62445 154245 0 0 $X=62305 $Y=153535
X166 2 VIA1_C_CDNS_724652447324 $T=63145 139255 0 0 $X=63005 $Y=138545
X167 2 VIA1_C_CDNS_724652447324 $T=63145 154245 0 0 $X=63005 $Y=153535
X168 2 VIA1_C_CDNS_724652447324 $T=68685 139255 0 0 $X=68545 $Y=138545
X169 2 VIA1_C_CDNS_724652447324 $T=68685 154245 0 0 $X=68545 $Y=153535
X170 2 VIA1_C_CDNS_724652447324 $T=79370 139430 0 0 $X=79230 $Y=138720
X171 4 VIA1_C_CDNS_724652447324 $T=81420 159580 0 0 $X=81280 $Y=158870
X172 7 VIA1_C_CDNS_724652447324 $T=82460 157800 0 0 $X=82320 $Y=157090
X173 4 VIA1_C_CDNS_724652447324 $T=83160 159580 0 0 $X=83020 $Y=158870
X174 8 VIA1_C_CDNS_724652447324 $T=84200 156020 0 0 $X=84060 $Y=155310
X175 8 VIA1_C_CDNS_724652447324 $T=84910 137650 0 0 $X=84770 $Y=136940
X176 2 VIA1_C_CDNS_724652447324 $T=85610 139430 0 0 $X=85470 $Y=138720
X177 7 VIA1_C_CDNS_724652447324 $T=91150 135870 0 0 $X=91010 $Y=135160
X178 9 VIA1_C_CDNS_724652447325 $T=81940 167700 0 0 $X=81020 $Y=167510
X179 7 VIA1_C_CDNS_724652447325 $T=82140 146820 0 0 $X=81220 $Y=146630
X180 10 VIA1_C_CDNS_724652447325 $T=83680 166920 0 0 $X=82760 $Y=166730
X181 7 VIA1_C_CDNS_724652447325 $T=88380 146820 0 0 $X=87460 $Y=146630
X182 2 VIA1_C_CDNS_724652447326 $T=15625 14715 0 0 $X=15485 $Y=13225
X183 2 VIA1_C_CDNS_724652447326 $T=15625 72555 0 0 $X=15485 $Y=71065
X184 6 VIA1_C_CDNS_724652447326 $T=40895 69275 0 0 $X=40755 $Y=67785
X185 6 VIA1_C_CDNS_724652447326 $T=40895 127115 0 0 $X=40755 $Y=125625
X186 2 VIA1_C_CDNS_724652447326 $T=66165 14715 0 0 $X=66025 $Y=13225
X187 2 VIA1_C_CDNS_724652447326 $T=66165 72555 0 0 $X=66025 $Y=71065
X188 2 VIA1_C_CDNS_724652447326 $T=68625 14715 0 0 $X=68485 $Y=13225
X189 2 VIA1_C_CDNS_724652447326 $T=68625 72555 0 0 $X=68485 $Y=71065
X190 6 VIA1_C_CDNS_724652447326 $T=93895 69275 0 0 $X=93755 $Y=67785
X191 6 VIA1_C_CDNS_724652447326 $T=93895 127115 0 0 $X=93755 $Y=125625
X192 2 VIA1_C_CDNS_724652447326 $T=119165 14715 0 0 $X=119025 $Y=13225
X193 2 VIA1_C_CDNS_724652447326 $T=119165 72555 0 0 $X=119025 $Y=71065
X194 2 VIA1_C_CDNS_724652447326 $T=121625 14715 0 0 $X=121485 $Y=13225
X195 2 VIA1_C_CDNS_724652447326 $T=121625 72555 0 0 $X=121485 $Y=71065
X196 6 VIA1_C_CDNS_724652447326 $T=146895 69275 0 0 $X=146755 $Y=67785
X197 6 VIA1_C_CDNS_724652447326 $T=146895 127115 0 0 $X=146755 $Y=125625
X198 2 VIA1_C_CDNS_724652447326 $T=172165 14715 0 0 $X=172025 $Y=13225
X199 2 VIA1_C_CDNS_724652447326 $T=172165 72555 0 0 $X=172025 $Y=71065
X200 2 VIA1_C_CDNS_724652447326 $T=174625 14715 0 0 $X=174485 $Y=13225
X201 2 VIA1_C_CDNS_724652447326 $T=174625 72555 0 0 $X=174485 $Y=71065
X202 6 VIA1_C_CDNS_724652447326 $T=199895 69275 0 0 $X=199755 $Y=67785
X203 6 VIA1_C_CDNS_724652447326 $T=199895 127115 0 0 $X=199755 $Y=125625
X204 2 VIA1_C_CDNS_724652447326 $T=225165 14715 0 0 $X=225025 $Y=13225
X205 2 VIA1_C_CDNS_724652447326 $T=225165 72555 0 0 $X=225025 $Y=71065
X206 2 VIA1_C_CDNS_724652447326 $T=227625 14715 0 0 $X=227485 $Y=13225
X207 2 VIA1_C_CDNS_724652447326 $T=227625 72555 0 0 $X=227485 $Y=71065
X208 6 VIA1_C_CDNS_724652447326 $T=252895 69275 0 0 $X=252755 $Y=67785
X209 6 VIA1_C_CDNS_724652447326 $T=252895 127115 0 0 $X=252755 $Y=125625
X210 2 VIA1_C_CDNS_724652447326 $T=278165 14715 0 0 $X=278025 $Y=13225
X211 2 VIA1_C_CDNS_724652447326 $T=278165 72555 0 0 $X=278025 $Y=71065
X212 6 2 VIA2_C_CDNS_724652447327 $T=10035 69275 0 0 $X=8545 $Y=67835
X213 6 2 VIA2_C_CDNS_724652447327 $T=10035 127115 0 0 $X=8545 $Y=125675
X214 2 2 VIA2_C_CDNS_724652447327 $T=13315 14715 0 0 $X=11825 $Y=13275
X215 2 2 VIA2_C_CDNS_724652447327 $T=13315 72555 0 0 $X=11825 $Y=71115
X216 2 2 VIA2_C_CDNS_724652447327 $T=280475 14715 0 0 $X=278985 $Y=13275
X217 2 2 VIA2_C_CDNS_724652447327 $T=280475 72555 0 0 $X=278985 $Y=71115
X218 6 2 VIA2_C_CDNS_724652447327 $T=283755 69275 0 0 $X=282265 $Y=67835
X219 6 2 VIA2_C_CDNS_724652447327 $T=283755 127115 0 0 $X=282265 $Y=125675
X220 3 VIA1_C_CDNS_7246524473210 $T=102805 160660 0 0 $X=100755 $Y=160170
X221 10 VIA1_C_CDNS_7246524473210 $T=124160 136175 0 0 $X=122110 $Y=135685
X222 3 VIA1_C_CDNS_7246524473210 $T=290340 136245 0 0 $X=288290 $Y=135755
X223 3 2 6 11 STE_3VX4 $T=97905 155845 0 0 $X=97475 $Y=155205
X224 2 8 6 ne3_CDNS_724652447320 $T=93475 156435 0 0 $X=92675 $Y=155905
X225 2 7 8 ne3_CDNS_724652447322 $T=79640 140720 0 0 $X=78840 $Y=140320
X226 2 7 7 ne3_CDNS_724652447322 $T=85880 140720 0 0 $X=85080 $Y=140320
X227 4 9 7 3 2 pe3_CDNS_724652447323 $T=81690 161500 0 0 $X=80180 $Y=160470
X228 4 10 8 3 2 pe3_CDNS_724652447323 $T=83430 161500 0 0 $X=81920 $Y=160470
X229 2 10 rpp1k1_3_CDNS_724652447324 $T=301000 19305 1 90 $X=300780 $Y=14145
X230 10 3 2 rpp1k1_3_CDNS_724652447327 $T=292340 141005 0 90 $X=121980 $Y=135845
X231 3 3 3 5 4 2 MASCO__A1 $T=25645 178655 0 0 $X=25645 $Y=178655
X232 3 3 3 5 5 2 MASCO__A1 $T=25645 196715 0 0 $X=25645 $Y=196715
X233 3 3 3 5 4 2 MASCO__A1 $T=25645 214775 0 0 $X=25645 $Y=214775
X234 3 5 5 5 4 2 MASCO__A1 $T=38125 178655 0 0 $X=38125 $Y=178655
X235 3 5 4 5 6 2 MASCO__A1 $T=38125 196715 0 0 $X=38125 $Y=196715
X236 3 5 5 5 4 2 MASCO__A1 $T=38125 214775 0 0 $X=38125 $Y=214775
X237 3 5 5 5 4 2 MASCO__A1 $T=50605 178655 0 0 $X=50605 $Y=178655
X238 3 5 4 5 5 2 MASCO__A1 $T=50605 196715 0 0 $X=50605 $Y=196715
X239 3 5 5 5 4 2 MASCO__A1 $T=50605 214775 0 0 $X=50605 $Y=214775
X240 3 5 5 5 4 2 MASCO__A1 $T=63085 178655 0 0 $X=63085 $Y=178655
X241 3 5 6 5 5 2 MASCO__A1 $T=63085 196715 0 0 $X=63085 $Y=196715
X242 3 5 5 5 4 2 MASCO__A1 $T=63085 214775 0 0 $X=63085 $Y=214775
X243 3 5 5 3 3 2 MASCO__A1 $T=75565 178655 0 0 $X=75565 $Y=178655
X244 3 3 3 3 3 2 MASCO__A1 $T=75565 196715 0 0 $X=75565 $Y=196715
X245 3 3 3 3 3 2 MASCO__A1 $T=75565 214775 0 0 $X=75565 $Y=214775
X246 2 2 1 1 MASCO__A2 $T=18935 140345 0 0 $X=18935 $Y=140345
X247 2 2 1 1 MASCO__A2 $T=18935 155315 0 0 $X=18935 $Y=155315
X248 2 1 5 1 MASCO__A2 $T=31415 140345 0 0 $X=31415 $Y=140345
X249 2 1 1 1 MASCO__A2 $T=31415 155315 0 0 $X=31415 $Y=155315
X250 2 1 1 1 MASCO__A2 $T=43895 140345 0 0 $X=43895 $Y=140345
X251 2 1 1 1 MASCO__A2 $T=43895 155315 0 0 $X=43895 $Y=155315
X252 2 1 2 2 MASCO__A2 $T=56375 140345 0 0 $X=56375 $Y=140345
X253 2 2 2 2 MASCO__A2 $T=56375 155315 0 0 $X=56375 $Y=155315
X254 6 2 2 MOSVC3 w=5e-05 l=5e-05 $X=15895 $Y=16925 $dt=2
X255 6 2 2 MOSVC3 w=5e-05 l=5e-05 $X=15895 $Y=74765 $dt=2
X256 6 2 2 MOSVC3 w=5e-05 l=5e-05 $X=68895 $Y=16925 $dt=2
X257 6 2 2 MOSVC3 w=5e-05 l=5e-05 $X=68895 $Y=74765 $dt=2
X258 6 2 2 MOSVC3 w=5e-05 l=5e-05 $X=121895 $Y=16925 $dt=2
X259 6 2 2 MOSVC3 w=5e-05 l=5e-05 $X=121895 $Y=74765 $dt=2
X260 6 2 2 MOSVC3 w=5e-05 l=5e-05 $X=174895 $Y=16925 $dt=2
X261 6 2 2 MOSVC3 w=5e-05 l=5e-05 $X=174895 $Y=74765 $dt=2
X262 6 2 2 MOSVC3 w=5e-05 l=5e-05 $X=227895 $Y=16925 $dt=2
X263 6 2 2 MOSVC3 w=5e-05 l=5e-05 $X=227895 $Y=74765 $dt=2
D10 2 3 p_dnw AREA=2.52272e-09 PJ=0.00028212 perimeter=0.00028212 $X=17665 $Y=173815 $dt=3
D11 2 3 p_dnw AREA=8.09228e-11 PJ=4.5e-05 perimeter=4.5e-05 $X=79040 $Y=154130 $dt=3
D12 2 2 p_dnw3 AREA=1.24376e-10 PJ=0.00020492 perimeter=0.00020492 $X=15095 $Y=16495 $dt=4
D13 2 2 p_dnw3 AREA=1.24376e-10 PJ=0.00020492 perimeter=0.00020492 $X=15095 $Y=74335 $dt=4
D14 2 3 p_dnw3 AREA=7.74011e-10 PJ=0 perimeter=0 $X=25645 $Y=178655 $dt=4
D15 2 3 p_dnw3 AREA=7.74011e-10 PJ=0 perimeter=0 $X=25645 $Y=196715 $dt=4
D16 2 3 p_dnw3 AREA=7.74011e-10 PJ=0 perimeter=0 $X=25645 $Y=214775 $dt=4
D17 2 2 p_dnw3 AREA=1.24376e-10 PJ=0.00020492 perimeter=0.00020492 $X=68095 $Y=16495 $dt=4
D18 2 2 p_dnw3 AREA=1.24376e-10 PJ=0.00020492 perimeter=0.00020492 $X=68095 $Y=74335 $dt=4
D19 2 3 p_dnw3 AREA=3.18756e-11 PJ=0 perimeter=0 $X=80180 $Y=160470 $dt=4
D20 2 2 p_dnw3 AREA=1.24376e-10 PJ=0.00020492 perimeter=0.00020492 $X=121095 $Y=16495 $dt=4
D21 2 2 p_dnw3 AREA=1.24376e-10 PJ=0.00020492 perimeter=0.00020492 $X=121095 $Y=74335 $dt=4
D22 2 2 p_dnw3 AREA=1.24376e-10 PJ=0.00020492 perimeter=0.00020492 $X=174095 $Y=16495 $dt=4
D23 2 2 p_dnw3 AREA=1.24376e-10 PJ=0.00020492 perimeter=0.00020492 $X=174095 $Y=74335 $dt=4
D24 2 2 p_dnw3 AREA=1.24376e-10 PJ=0.00020492 perimeter=0.00020492 $X=227095 $Y=16495 $dt=4
D25 2 2 p_dnw3 AREA=1.24376e-10 PJ=0.00020492 perimeter=0.00020492 $X=227095 $Y=74335 $dt=4
.ends por2
