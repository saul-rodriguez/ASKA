************************************************************************
* auCdl Netlist:
* 
* Library Name:  ASKA_PULSE_GENERATOR
* Top Cell Name: pulse_generator
* View Name:     schematic
* Netlisted on:  Aug 26 08:46:57 2024
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.LDD
*.SCALE METER
.PARAM



************************************************************************
* Library Name: ASKA_CURRENT_SOURCE
* Cell Name:    current_source_gm_10_en_r
* View Name:    schematic
************************************************************************

.SUBCKT current_source_gm_10_en_r BIAS EN FB GNDA GNDHV IN OUT PACTIVE VDD3A 
+ VDDHV VSUBHV
*.PININFO BIAS:B EN:B FB:B GNDA:B GNDHV:B IN:B OUT:B PACTIVE:B VDD3A:B VDDHV:B 
*.PININFO VSUBHV:B
XC0 VDD3A GNDA GNDA / mosvc3 W=20u L=30u M=4.0 par1=4.0
MM30 VDD3A VDD3A VDD3A VDD3A PE3 W=10u L=5u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM26 net16 EN VDD3A VDD3A PE3 W=3u L=300n M=2.0 AD=2.88e-12 AS=2.88e-12 
+ PD=1.296e-05 PS=1.296e-05 NRD=0.045 NRS=0.045
MM35 net13 PACTIVE VDD3A VDD3A PE3 W=3u L=300n M=2.0 AD=2.88e-12 AS=2.88e-12 
+ PD=1.296e-05 PS=1.296e-05 NRD=0.045 NRS=0.045
MM23 net15 net15 VDD3A VDD3A PE3 W=10u L=1u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM29 VDD3A VDD3A VDD3A VDD3A PE3 W=10u L=5u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM11 net10 net4 VDD3A VDD3A PE3 W=10u L=5u M=2.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM9 net6 net4 VDD3A VDD3A PE3 W=10u L=5u M=2.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM10 net8 net4 VDD3A VDD3A PE3 W=10u L=5u M=20.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM20 VB net15 VDD3A VDD3A PE3 W=10u L=1u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM5 net9 net10 net8 VDD3A PE3 W=10u L=5u M=14.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM3 net7 net6 net8 VDD3A PE3 W=10u L=5u M=14.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM12 net4 net4 VDD3A VDD3A PE3 W=10u L=5u M=2.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM8 GNDA IN net6 net6 PE3 W=10u L=5u M=18.0 AD=2.93333e-12 AS=2.93333e-12 
+ PD=1.16978e-05 PS=1.16978e-05 NRD=0.027 NRS=0.027
MM7 GNDA net1 net10 net10 PE3 W=10u L=5u M=18.0 AD=2.93333e-12 AS=2.93333e-12 
+ PD=1.16978e-05 PS=1.16978e-05 NRD=0.027 NRS=0.027
MM25 net16 EN GNDA GNDA NE3 W=2u L=350.0n M=1.0 AD=9.6e-13 AS=9.6e-13 
+ PD=4.96e-06 PS=4.96e-06 NRD=0.135 NRS=0.135
MM24 net12 net16 GNDA GNDA NE3 W=5u L=350.0n M=4.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM34 net13 PACTIVE GNDA GNDA NE3 W=2u L=350.0n M=1.0 AD=9.6e-13 AS=9.6e-13 
+ PD=4.96e-06 PS=4.96e-06 NRD=0.135 NRS=0.135
MM32 net9 net13 GNDA GNDA NE3 W=5u L=350.0n M=4.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM22 net15 BIAS net14 GNDA NE3 W=10u L=10u M=2.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM21 net14 net12 GNDA GNDA NE3 W=10u L=10u M=2.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM19 net4 BIAS net5 GNDA NE3 W=10u L=10u M=2.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM18 BIAS BIAS net12 GNDA NE3 W=10u L=10u M=2.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM27 GNDA GNDA GNDA GNDA NE3 W=10u L=10u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM6 VB net9 GNDA GNDA NE3 W=5u L=500n M=4.0 AD=1.35e-12 AS=1.875e-12 
+ PD=5.54e-06 PS=8.25e-06 NRD=0.054 NRS=0.054
MM4 net7 net7 GNDA GNDA NE3 W=5u L=1u M=2.0 AD=2.4e-12 AS=2.4e-12 PD=1.096e-05 
+ PS=1.096e-05 NRD=0.054 NRS=0.054
MM2 net9 net7 GNDA GNDA NE3 W=5u L=1u M=2.0 AD=2.4e-12 AS=2.4e-12 PD=1.096e-05 
+ PS=1.096e-05 NRD=0.054 NRS=0.054
MM13 net5 net12 GNDA GNDA NE3 W=10u L=10u M=2.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM14 net12 net12 GNDA GNDA NE3 W=10u L=10u M=2.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM0 OUT VA FB VSUBHV NEDIA W=100.0000u L=1.25u M=8.0 $LDD[NEDIA]
MM1 VA VB GNDHV VSUBHV NEDIA W=50u L=1.25u M=1.0 $LDD[NEDIA]
RR1 VSUBHV GNDA 5.0 $[S_RES]
CC1 net9 net11 $[CMM5T] area=8.4e-10 perimeter=116.000000u M=7
RR7 GNDHV OUT 1.00618M $SUB=VSUBHV $[RPP1K1_3] $W=2u $L=2.04358m M=1
RR4 FB net1 5031.08 $SUB=GNDA $[RPP1K1_3] $W=2u $L=10u M=9
RR2 VA VDDHV 99.9954K $SUB=VSUBHV $[RPP1K1_3] $W=4u $L=411.22u M=1
RR3 GNDHV VA 25.0012K $SUB=VSUBHV $[RPP1K1_3] $W=4u $L=102.65u M=1
RR0 net11 VB 39.9966K $SUB=VDD3A $[RPP1K1_3] $W=4u $L=164.35u M=1
.ENDS

************************************************************************
* Library Name: ASKA_DAC6B
* Cell Name:    dac6b_amp_n2
* View Name:    schematic
************************************************************************

.SUBCKT dac6b_amp_n2 BIAS D0 D1 D2 D3 D4 D5 ENABLE GNDA VDDA VOUT VREF
*.PININFO BIAS:B D0:B D1:B D2:B D3:B D4:B D5:B ENABLE:B GNDA:B VDDA:B VOUT:B 
*.PININFO VREF:B
MM43 VDDA VDDA VDDA VDDA PE3 W=2u L=10u M=30.0 AD=9.6e-13 AS=9.6e-13 
+ PD=4.96e-06 PS=4.96e-06 NRD=0.135 NRS=0.135
MM42 VDDA VDDA VDDA VDDA PE3 W=10u L=10u M=17.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM36 VDDA VDDA VDDA VDDA PE3 W=10u L=10u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM35 EN ENABLE VDDA VDDA PE3 W=6u L=300n M=1.0 AD=2.88e-12 AS=2.88e-12 
+ PD=1.296e-05 PS=1.296e-05 NRD=0.045 NRS=0.045
MM31 GNDA GNDA net34 net34 PE3 W=10u L=20u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM30 net34 net34 net30 net30 PE3 W=10u L=20u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM29 net30 net30 net10 net10 PE3 W=10u L=20u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM28 net8 net8 VDDA VDDA PE3 W=10u L=10u M=2.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM27 net10 net8 VDDA VDDA PE3 W=10u L=10u M=2.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM23 net12 net12 VDDA VDDA PE3 W=10u L=10u M=8.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM21 net14 net30 net19 VDDA PE3 W=10u L=1u M=10.0 AD=2.7e-12 AS=3.12e-12 
+ PD=1.054e-05 PS=1.2624e-05 NRD=0.027 NRS=0.027
MM20 GNDA D5 net5 VDDA PE3 W=10u L=350.0n M=2.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM19 GNDA D4 net4 VDDA PE3 W=10u L=350.0n M=2.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM18 GNDA D3 net3 VDDA PE3 W=10u L=350.0n M=2.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM17 GNDA D2 net2 VDDA PE3 W=10u L=350.0n M=2.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM16 GNDA D1 net1 VDDA PE3 W=10u L=350.0n M=2.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM15 GNDA D0 net6 VDDA PE3 W=10u L=350.0n M=2.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM14 net19 net7 VDDA VDDA PE3 W=10u L=10u M=10.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM22 net7 net12 VDDA VDDA PE3 W=10u L=10u M=8.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM11 VOUT net30 net5 VDDA PE3 W=10u L=1u M=32.0 AD=2.7e-12 AS=2.83125e-12 
+ PD=1.054e-05 PS=1.11913e-05 NRD=0.027 NRS=0.027
MM10 VOUT net30 net4 VDDA PE3 W=10u L=1u M=16.0 AD=2.7e-12 AS=2.9625e-12 
+ PD=1.054e-05 PS=1.18425e-05 NRD=0.027 NRS=0.027
MM9 VOUT net30 net3 VDDA PE3 W=10u L=1u M=8.0 AD=2.7e-12 AS=3.225e-12 
+ PD=1.054e-05 PS=1.3145e-05 NRD=0.027 NRS=0.027
MM8 VOUT net30 net2 VDDA PE3 W=10u L=1u M=4.0 AD=2.7e-12 AS=3.75e-12 
+ PD=1.054e-05 PS=1.575e-05 NRD=0.027 NRS=0.027
MM7 VOUT net30 net1 VDDA PE3 W=10u L=1u M=2.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM6 VOUT net30 net6 VDDA PE3 W=10u L=1u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM5 net5 net7 VDDA VDDA PE3 W=10u L=10u M=32.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM4 net4 net7 VDDA VDDA PE3 W=10u L=10u M=16.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM3 net3 net7 VDDA VDDA PE3 W=10u L=10u M=8.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM2 net2 net7 VDDA VDDA PE3 W=10u L=10u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM1 net1 net7 VDDA VDDA PE3 W=10u L=10u M=2.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM0 net6 net7 VDDA VDDA PE3 W=10u L=10u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
RR1 GNDA net14 200.001K $SUB=GNDA $[RPP1K1_3] $W=4u $L=822.7u M=1
RR0 GNDA VOUT 52.7974K $SUB=GNDA $[RPP1K1_3] $W=4u $L=217.02u M=1
XM41 A A A A VDDA GNDA / ne3i_6 W=10u L=2u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ NRD=0.027 NRS=0.027 PD=2.096e-05 PS=2.096e-05 par1=4.0
XM12 net7 VREF A A VDDA GNDA / ne3i_6 W=10u L=2u M=16.0 AD=4.8e-12 AS=4.8e-12 
+ NRD=0.027 NRS=0.027 PD=2.096e-05 PS=2.096e-05 par1=16.0
XM24 net12 net14 A A VDDA GNDA / ne3i_6 W=10u L=2u M=16.0 AD=4.8e-12 
+ AS=4.8e-12 NRD=0.027 NRS=0.027 PD=2.096e-05 PS=2.096e-05 par1=16.0
MM40 GNDA GNDA GNDA GNDA NE3 W=10u L=2u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM38 A BIAS net15 GNDA NE3 W=10u L=2u M=8.0 AD=2.7e-12 AS=3.225e-12 
+ PD=1.054e-05 PS=1.3145e-05 NRD=0.027 NRS=0.027
MM37 net8 BIAS net13 GNDA NE3 W=10u L=2u M=8.0 AD=2.7e-12 AS=3.225e-12 
+ PD=1.054e-05 PS=1.3145e-05 NRD=0.027 NRS=0.027
MM39 BIAS BIAS net9 GNDA NE3 W=10u L=2u M=8.0 AD=2.7e-12 AS=3.225e-12 
+ PD=1.054e-05 PS=1.3145e-05 NRD=0.027 NRS=0.027
MM34 EN ENABLE GNDA GNDA NE3 W=2u L=350.0n M=1.0 AD=9.6e-13 AS=9.6e-13 
+ PD=4.96e-06 PS=4.96e-06 NRD=0.135 NRS=0.135
MM33 net9 EN GNDA GNDA NE3 W=10u L=350.0n M=4.0 AD=2.7e-12 AS=3.75e-12 
+ PD=1.054e-05 PS=1.575e-05 NRD=0.027 NRS=0.027
MM26 net13 net9 GNDA GNDA NE3 W=10u L=2u M=8.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM13 net9 net9 GNDA GNDA NE3 W=10u L=2u M=8.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM25 net15 net9 GNDA GNDA NE3 W=10u L=2u M=8.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM32 VOUT EN GNDA GNDA NE3 W=10u L=350.0n M=4.0 AD=2.7e-12 AS=3.75e-12 
+ PD=1.054e-05 PS=1.575e-05 NRD=0.027 NRS=0.027
.ENDS

************************************************************************
* Library Name: ASKA_PULSE_GENERATOR
* Cell Name:    pulse_generator
* View Name:    schematic
************************************************************************

.SUBCKT pulse_generator BIAS1 BIAS2 CUR_OUT D<5> D<4> D<3> D<2> D<1> D<0> 
+ ENABLE EXT_FB_RES GNDA GNDHV PULSE_ACTIVE VDD3A VDDHV VREF VSUBHV
*.PININFO BIAS1:B BIAS2:B CUR_OUT:B D<5>:B D<4>:B D<3>:B D<2>:B D<1>:B D<0>:B 
*.PININFO ENABLE:B EXT_FB_RES:B GNDA:B GNDHV:B PULSE_ACTIVE:B VDD3A:B VDDHV:B 
*.PININFO VREF:B VSUBHV:B
XC1 VDD3A GNDA GNDA / mosvc3 W=20u L=20u M=8.0 par1=8.0
XC0 VDD3A GNDA GNDA / mosvc3 W=25.0u L=20u M=4.0 par1=4.0
XI1 BIAS2 ENABLE EXT_FB_RES GNDA GNDHV VDAC CUR_OUT PULSE_ACTIVE VDD3A VDDHV 
+ VSUBHV / current_source_gm_10_en_r
XI0 BIAS1 D<0> D<1> D<2> D<3> D<4> D<5> ENABLE GNDA VDD3A VDAC VREF / 
+ dac6b_amp_n2
.ENDS


.SUBCKT ne3i_6 D G S B NW SB 
*.PININFO  D:B G:B S:B B:B NW:B SB:B
.ENDS

.SUBCKT mosvc3 G NW SB 
*.PININFO  G:B NW:B SB:B
.ENDS
