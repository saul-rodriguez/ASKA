* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : current_source_gm_10_en_r                    *
* Netlisted  : Tue Aug 13 03:37:13 2024                     *
* PVS Version: 23.10-p043 Mon Oct 2 18:09:08 PDT 2023      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 LDDN(nedia) nedia2_d dnwtrm(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 1 MN(ne3) nem ndiff(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 2 MP(pe3) pem pdiff(D) p1trm(G) pdiff(S) nwtrm(B)
*.DEVTMPLT 3 MOSVC3() mosvcm p1trm(G) nwtrm(NW) bulk(SB)
*.DEVTMPLT 4 R(s_res) s_res bulk(POS) bulk(NEG)
*.DEVTMPLT 5 D(p_dnw) p_dnw bulk(POS) nwtrm(NEG)
*.DEVTMPLT 6 D(p_dnw3) p_dnwm bulk(POS) nwtrm(NEG)
*.DEVTMPLT 7 R(rpp1k1_3) rpp1k1_s p1trm(POS) p1trm(NEG) bulk(SUB)
*.DEVTMPLT 8 R(rpp1k1_3) rpp1k1_n p1trm(POS) p1trm(NEG) nwtrm(SUB)
*.DEVTMPLT 9 C(cmm5t) cmim capm(POS) m4trm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_723534627840                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_723534627840 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_723534627840

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_723534627841                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_723534627841 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_723534627841

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_723534627842                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_723534627842 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_723534627842

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_723534627843                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_723534627843 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_723534627843

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_723534627844                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_723534627844 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_723534627844

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_723534627845                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_723534627845 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_723534627845

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_723534627846                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_723534627846 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_723534627846

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_723534627847                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_723534627847 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_723534627847

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_723534627848                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_723534627848 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_723534627848

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_723534627849                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_723534627849 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_723534627849

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7235346278410                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7235346278410 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7235346278410

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ND_C_CDNS_7235346278411                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ND_C_CDNS_7235346278411 1 2
** N=2 EP=2 FDC=0
.ends ND_C_CDNS_7235346278411

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7235346278412                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7235346278412 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7235346278412

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7235346278413                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7235346278413 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7235346278413

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7235346278414                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7235346278414 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7235346278414

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7235346278416                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7235346278416 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7235346278416

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7235346278417                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7235346278417 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7235346278417

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7235346278418                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7235346278418 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7235346278418

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7235346278419                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7235346278419 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7235346278419

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7235346278420                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7235346278420 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7235346278420

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7235346278422                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7235346278422 1 2
** N=2 EP=2 FDC=0
.ends VIA2_C_CDNS_7235346278422

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7235346278423                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7235346278423 1 2
** N=2 EP=2 FDC=0
.ends VIA1_C_CDNS_7235346278423

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_7235346278432                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_7235346278432 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_7235346278432

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7235346278438                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7235346278438 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7235346278438

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7235346278440                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7235346278440 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7235346278440

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7235346278444                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7235346278444 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7235346278444

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7235346278453                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7235346278453 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7235346278453

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_723534627840                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_723534627840 1 2 3
** N=3 EP=3 FDC=4
M0 3 2 1 1 ne3 L=5e-07 W=5e-06 AD=1.35e-12 AS=2.4e-12 PD=5.54e-06 PS=1.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 1 ne3 L=5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=1040 $Y=0 $dt=1
M2 3 2 1 1 ne3 L=5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=2080 $Y=0 $dt=1
M3 1 2 3 1 ne3 L=5e-07 W=5e-06 AD=2.4e-12 AS=1.35e-12 PD=1.096e-05 PS=5.54e-06 $X=3120 $Y=0 $dt=1
.ends ne3_CDNS_723534627840

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nedia_CDNS_723534627841                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nedia_CDNS_723534627841 1 2 3 4
** N=4 EP=4 FDC=1
X0 2 4 3 1 LDDN w=5e-05 l=1.25e-06 adio=1.08602e-09 pdio=0.00013535 extlay=1 $[nedia] $X=-680 $Y=-4850 $dt=0
.ends nedia_CDNS_723534627841

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_723534627842                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_723534627842 1 2 3
** N=3 EP=3 FDC=4
M0 3 2 1 1 ne3 L=3.5e-07 W=5e-06 AD=1.35e-12 AS=2.4e-12 PD=5.54e-06 PS=1.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 1 ne3 L=3.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=890 $Y=0 $dt=1
M2 3 2 1 1 ne3 L=3.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=1780 $Y=0 $dt=1
M3 1 2 3 1 ne3 L=3.5e-07 W=5e-06 AD=2.4e-12 AS=1.35e-12 PD=1.096e-05 PS=5.54e-06 $X=2670 $Y=0 $dt=1
.ends ne3_CDNS_723534627842

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_723534627843                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_723534627843 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.00010265 W=4e-06 $[rpp1k1_3] $SUB=3 $X=0 $Y=0 $dt=7
.ends rpp1k1_3_CDNS_723534627843

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nedia_CDNS_723534627844                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nedia_CDNS_723534627844 1 2 3 4
** N=4 EP=4 FDC=8
X0 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=-680 $Y=-4850 $dt=0
X1 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=11220 $Y=-4850 $dt=0
X2 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=23120 $Y=-4850 $dt=0
X3 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=35020 $Y=-4850 $dt=0
X4 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=46920 $Y=-4850 $dt=0
X5 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=58820 $Y=-4850 $dt=0
X6 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=70720 $Y=-4850 $dt=0
X7 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=82620 $Y=-4850 $dt=0
.ends nedia_CDNS_723534627844

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_723534627845                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_723534627845 1 2 3 4
** N=4 EP=4 FDC=2
M0 3 2 1 4 ne3 L=1e-05 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 ne3 L=1e-05 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=10540 $Y=0 $dt=1
.ends ne3_CDNS_723534627845

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_723534627846                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_723534627846 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
M0 3 2 1 1 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
.ends pe3_CDNS_723534627846

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_723534627847                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_723534627847 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=2
M0 3 2 1 1 pe3 L=3e-07 W=3e-06 AD=8.1e-13 AS=1.44e-12 PD=3.54e-06 PS=6.96e-06 $X=0 $Y=0 $dt=2
M1 1 2 3 1 pe3 L=3e-07 W=3e-06 AD=1.44e-12 AS=8.1e-13 PD=6.96e-06 PS=3.54e-06 $X=840 $Y=0 $dt=2
.ends pe3_CDNS_723534627847

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_723534627848                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_723534627848 1 2 3
** N=3 EP=3 FDC=1
R0 1 2 L=0.00204354 W=2e-06 $[rpp1k1_3] $SUB=3 $X=-2220 $Y=0 $dt=7
.ends rpp1k1_3_CDNS_723534627848

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7235346278411                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7235346278411 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=1
M0 3 2 1 4 pe3 L=5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
.ends pe3_CDNS_7235346278411

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7235346278412                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7235346278412 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=1e-05 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends ne3_CDNS_7235346278412

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7235346278413                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7235346278413 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=1e-06 W=5e-06 AD=2.4e-12 AS=2.4e-12 PD=1.096e-05 PS=1.096e-05 $X=0 $Y=0 $dt=1
.ends ne3_CDNS_7235346278413

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7235346278414                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7235346278414 1 2 3
*.DEVICECLIMB
** N=3 EP=3 FDC=9
M0 3 2 1 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
M1 1 2 3 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=5540 $Y=0 $dt=2
M2 3 2 1 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=11080 $Y=0 $dt=2
M3 1 2 3 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=16620 $Y=0 $dt=2
M4 3 2 1 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=22160 $Y=0 $dt=2
M5 1 2 3 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=27700 $Y=0 $dt=2
M6 3 2 1 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=33240 $Y=0 $dt=2
M7 1 2 3 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=38780 $Y=0 $dt=2
M8 3 2 1 1 pe3 L=5e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=44320 $Y=0 $dt=2
.ends pe3_CDNS_7235346278414

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7235346278415                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7235346278415 1 2 3
** N=3 EP=3 FDC=1
R0 1 2 L=1e-05 W=2e-06 $[rpp1k1_3] $SUB=3 $X=0 $Y=0 $dt=7
.ends rpp1k1_3_CDNS_7235346278415

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7235346278416                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7235346278416 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
R0 2 1 L=0.00016435 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=8
.ends rpp1k1_3_CDNS_7235346278416

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7235346278417                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7235346278417 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.00041122 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=7
.ends rpp1k1_3_CDNS_7235346278417

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7235346278418                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7235346278418 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=3.5e-07 W=2e-06 AD=9.6e-13 AS=9.6e-13 PD=4.96e-06 PS=4.96e-06 $X=0 $Y=0 $dt=1
.ends ne3_CDNS_7235346278418

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7235346278443                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7235346278443 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7235346278443

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X1 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7235346278443 $T=660 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7235346278443 $T=660 1500 0 0 $X=0 $Y=1000
X2 1 VIATP_C_CDNS_7235346278443 $T=660 2500 0 0 $X=0 $Y=2000
X3 1 VIATP_C_CDNS_7235346278443 $T=660 3500 0 0 $X=0 $Y=3000
X4 1 VIATP_C_CDNS_7235346278443 $T=660 4500 0 0 $X=0 $Y=4000
.ends MASCO__X1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7235346278442                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7235346278442 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7235346278442

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X2 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7235346278442 $T=790 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7235346278442 $T=790 1500 0 0 $X=0 $Y=1000
X2 1 VIATP_C_CDNS_7235346278442 $T=790 2500 0 0 $X=0 $Y=2000
X3 1 VIATP_C_CDNS_7235346278442 $T=790 3500 0 0 $X=0 $Y=3000
X4 1 VIATP_C_CDNS_7235346278442 $T=790 4500 0 0 $X=0 $Y=4000
.ends MASCO__X2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7235346278439                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7235346278439 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7235346278439

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y6                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y6 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7235346278439 $T=500 530 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7235346278439 $T=1500 530 0 0 $X=1000 $Y=0
X2 1 VIATP_C_CDNS_7235346278439 $T=2500 530 0 0 $X=2000 $Y=0
X3 1 VIATP_C_CDNS_7235346278439 $T=3500 530 0 0 $X=3000 $Y=0
X4 1 VIATP_C_CDNS_7235346278439 $T=4500 530 0 0 $X=4000 $Y=0
X5 1 VIATP_C_CDNS_7235346278439 $T=5500 530 0 0 $X=5000 $Y=0
X6 1 VIATP_C_CDNS_7235346278439 $T=6500 530 0 0 $X=6000 $Y=0
X7 1 VIATP_C_CDNS_7235346278439 $T=7500 530 0 0 $X=7000 $Y=0
X8 1 VIATP_C_CDNS_7235346278439 $T=8500 530 0 0 $X=8000 $Y=0
X9 1 VIATP_C_CDNS_7235346278439 $T=9500 530 0 0 $X=9000 $Y=0
X10 1 VIATP_C_CDNS_7235346278439 $T=10500 530 0 0 $X=10000 $Y=0
.ends MASCO__Y6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7235346278441                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7235346278441 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7235346278441

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X5                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X5 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7235346278441 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7235346278441 $T=500 1500 0 0 $X=0 $Y=1000
X2 1 VIATP_C_CDNS_7235346278441 $T=500 2500 0 0 $X=0 $Y=2000
X3 1 VIATP_C_CDNS_7235346278441 $T=500 3500 0 0 $X=0 $Y=3000
X4 1 VIATP_C_CDNS_7235346278441 $T=500 4500 0 0 $X=0 $Y=4000
.ends MASCO__X5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y7                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y7 1
** N=1 EP=1 FDC=0
X0 1 MASCO__X5 $T=0 0 0 0 $X=0 $Y=0
X1 1 MASCO__X5 $T=2000 0 0 0 $X=2000 $Y=0
X2 1 MASCO__X5 $T=4000 0 0 0 $X=4000 $Y=0
X3 1 MASCO__X5 $T=6000 0 0 0 $X=6000 $Y=0
X4 1 MASCO__X5 $T=8000 0 0 0 $X=8000 $Y=0
X5 1 MASCO__X5 $T=10000 0 0 0 $X=10000 $Y=0
X6 1 MASCO__X5 $T=12000 0 0 0 $X=12000 $Y=0
X7 1 MASCO__X5 $T=14000 0 0 0 $X=14000 $Y=0
X8 1 MASCO__X5 $T=16000 0 0 0 $X=16000 $Y=0
.ends MASCO__Y7

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X4                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X4 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7235346278441 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7235346278441 $T=500 2500 0 0 $X=0 $Y=2000
X2 1 VIATP_C_CDNS_7235346278441 $T=500 4500 0 0 $X=0 $Y=4000
X3 1 VIATP_C_CDNS_7235346278441 $T=500 6500 0 0 $X=0 $Y=6000
X4 1 VIATP_C_CDNS_7235346278441 $T=500 8500 0 0 $X=0 $Y=8000
X5 1 VIATP_C_CDNS_7235346278441 $T=500 10500 0 0 $X=0 $Y=10000
X6 1 VIATP_C_CDNS_7235346278441 $T=500 12500 0 0 $X=0 $Y=12000
X7 1 VIATP_C_CDNS_7235346278441 $T=500 14500 0 0 $X=0 $Y=14000
X8 1 VIATP_C_CDNS_7235346278441 $T=500 16500 0 0 $X=0 $Y=16000
X9 1 VIATP_C_CDNS_7235346278441 $T=500 18500 0 0 $X=0 $Y=18000
X10 1 VIATP_C_CDNS_7235346278441 $T=500 20500 0 0 $X=0 $Y=20000
X11 1 VIATP_C_CDNS_7235346278441 $T=500 22500 0 0 $X=0 $Y=22000
.ends MASCO__X4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y8                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y8 1
** N=1 EP=1 FDC=0
X0 1 MASCO__X4 $T=0 0 0 0 $X=0 $Y=0
X1 1 MASCO__X4 $T=2000 0 0 0 $X=2000 $Y=0
X2 1 MASCO__X4 $T=4000 0 0 0 $X=4000 $Y=0
X3 1 MASCO__X4 $T=6000 0 0 0 $X=6000 $Y=0
X4 1 MASCO__X4 $T=8000 0 0 0 $X=8000 $Y=0
X5 1 MASCO__X4 $T=10000 0 0 0 $X=10000 $Y=0
X6 1 MASCO__X4 $T=12000 0 0 0 $X=12000 $Y=0
.ends MASCO__Y8

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X3                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X3 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7235346278441 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7235346278441 $T=500 2500 0 0 $X=0 $Y=2000
X2 1 VIATP_C_CDNS_7235346278441 $T=500 4500 0 0 $X=0 $Y=4000
X3 1 VIATP_C_CDNS_7235346278441 $T=500 6500 0 0 $X=0 $Y=6000
X4 1 VIATP_C_CDNS_7235346278441 $T=500 8500 0 0 $X=0 $Y=8000
X5 1 VIATP_C_CDNS_7235346278441 $T=500 10500 0 0 $X=0 $Y=10000
X6 1 VIATP_C_CDNS_7235346278441 $T=500 12500 0 0 $X=0 $Y=12000
X7 1 VIATP_C_CDNS_7235346278441 $T=500 14500 0 0 $X=0 $Y=14000
X8 1 VIATP_C_CDNS_7235346278441 $T=500 16500 0 0 $X=0 $Y=16000
X9 1 VIATP_C_CDNS_7235346278441 $T=500 18500 0 0 $X=0 $Y=18000
X10 1 VIATP_C_CDNS_7235346278441 $T=500 20500 0 0 $X=0 $Y=20000
.ends MASCO__X3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y9                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y9 1
** N=1 EP=1 FDC=0
X0 1 MASCO__X3 $T=0 0 0 0 $X=0 $Y=0
X1 1 MASCO__X3 $T=2000 0 0 0 $X=2000 $Y=0
X2 1 MASCO__X3 $T=4000 0 0 0 $X=4000 $Y=0
X3 1 MASCO__X3 $T=6000 0 0 0 $X=6000 $Y=0
X4 1 MASCO__X3 $T=8000 0 0 0 $X=8000 $Y=0
X5 1 MASCO__X3 $T=10000 0 0 0 $X=10000 $Y=0
X6 1 MASCO__X3 $T=12000 0 0 0 $X=12000 $Y=0
.ends MASCO__Y9

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: current_source_gm_10_en_r                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt current_source_gm_10_en_r 2 19 23 9 16 18 24 20 14 27
+ 25
** N=27 EP=11 FDC=198
X0 1 VIA1_C_CDNS_723534627840 $T=7790 61030 0 0 $X=7390 $Y=60320
X1 2 VIA1_C_CDNS_723534627840 $T=18330 62810 0 0 $X=17930 $Y=62100
X2 1 VIA1_C_CDNS_723534627840 $T=28870 61030 0 0 $X=28470 $Y=60320
X3 3 VIA1_C_CDNS_723534627840 $T=33575 62810 0 0 $X=33175 $Y=62100
X4 4 VIA1_C_CDNS_723534627840 $T=44115 61030 0 0 $X=43715 $Y=60320
X5 3 VIA1_C_CDNS_723534627840 $T=54655 62810 0 0 $X=54255 $Y=62100
X6 5 VIA1_C_CDNS_723534627840 $T=59300 62950 0 0 $X=58900 $Y=62240
X7 6 VIA1_C_CDNS_723534627840 $T=69840 61110 0 0 $X=69440 $Y=60400
X8 5 VIA1_C_CDNS_723534627840 $T=80380 62950 0 0 $X=79980 $Y=62240
X9 7 VIA1_C_CDNS_723534627840 $T=106545 17830 0 0 $X=106145 $Y=17120
X10 8 VIA1_C_CDNS_723534627840 $T=106545 45950 0 0 $X=106145 $Y=45240
X11 7 VIA1_C_CDNS_723534627840 $T=117625 17830 0 0 $X=117225 $Y=17120
X12 8 VIA1_C_CDNS_723534627840 $T=117625 45950 0 0 $X=117225 $Y=45240
X13 7 VIA1_C_CDNS_723534627840 $T=128705 17830 0 0 $X=128305 $Y=17120
X14 8 VIA1_C_CDNS_723534627840 $T=128705 45950 0 0 $X=128305 $Y=45240
X15 7 VIA1_C_CDNS_723534627840 $T=139785 17830 0 0 $X=139385 $Y=17120
X16 8 VIA1_C_CDNS_723534627840 $T=139785 45950 0 0 $X=139385 $Y=45240
X17 7 VIA1_C_CDNS_723534627840 $T=150865 17830 0 0 $X=150465 $Y=17120
X18 8 VIA1_C_CDNS_723534627840 $T=150865 45950 0 0 $X=150465 $Y=45240
X19 8 VIA1_C_CDNS_723534627840 $T=160825 16050 0 0 $X=160425 $Y=15340
X20 7 VIA1_C_CDNS_723534627840 $T=160825 47730 0 0 $X=160425 $Y=47020
X21 8 VIA1_C_CDNS_723534627840 $T=171905 16050 0 0 $X=171505 $Y=15340
X22 7 VIA1_C_CDNS_723534627840 $T=171905 47730 0 0 $X=171505 $Y=47020
X23 8 VIA1_C_CDNS_723534627840 $T=182985 16050 0 0 $X=182585 $Y=15340
X24 7 VIA1_C_CDNS_723534627840 $T=182985 47730 0 0 $X=182585 $Y=47020
X25 8 VIA1_C_CDNS_723534627840 $T=194065 16050 0 0 $X=193665 $Y=15340
X26 7 VIA1_C_CDNS_723534627840 $T=194065 47730 0 0 $X=193665 $Y=47020
X27 8 VIA1_C_CDNS_723534627840 $T=205145 16050 0 0 $X=204745 $Y=15340
X28 7 VIA1_C_CDNS_723534627840 $T=205145 47730 0 0 $X=204745 $Y=47020
X29 9 VIA1_C_CDNS_723534627841 $T=247850 19860 0 0 $X=247710 $Y=18890
X30 10 VIA1_C_CDNS_723534627841 $T=248890 17580 0 0 $X=248750 $Y=16610
X31 9 VIA1_C_CDNS_723534627841 $T=249930 19860 0 0 $X=249790 $Y=18890
X32 10 VIA1_C_CDNS_723534627841 $T=250970 17580 0 0 $X=250830 $Y=16610
X33 9 VIA1_C_CDNS_723534627841 $T=252010 19860 0 0 $X=251870 $Y=18890
X34 1 VIA1_C_CDNS_723534627842 $T=33660 31900 0 0 $X=33260 $Y=31710
X35 1 VIA1_C_CDNS_723534627842 $T=44900 31900 0 0 $X=44500 $Y=31710
X36 1 VIA1_C_CDNS_723534627842 $T=56140 31900 0 0 $X=55740 $Y=31710
X37 4 VIA1_C_CDNS_723534627842 $T=63465 83370 0 0 $X=63065 $Y=83180
X38 4 VIA1_C_CDNS_723534627842 $T=65705 83370 0 0 $X=65305 $Y=83180
X39 4 VIA1_C_CDNS_723534627842 $T=67945 83370 0 0 $X=67545 $Y=83180
X40 4 VIA1_C_CDNS_723534627842 $T=70185 83370 0 0 $X=69785 $Y=83180
X41 4 VIA1_C_CDNS_723534627842 $T=72425 83370 0 0 $X=72025 $Y=83180
X42 7 VIA1_C_CDNS_723534627842 $T=117900 81120 0 0 $X=117500 $Y=80930
X43 8 VIA1_C_CDNS_723534627842 $T=119550 81900 0 0 $X=119150 $Y=81710
X44 6 VIA1_C_CDNS_723534627842 $T=122400 137545 0 0 $X=122000 $Y=137355
X45 7 VIA1_C_CDNS_723534627842 $T=124680 81120 0 0 $X=124280 $Y=80930
X46 8 VIA1_C_CDNS_723534627842 $T=125360 81900 0 0 $X=124960 $Y=81710
X47 6 VIA1_C_CDNS_723534627842 $T=128640 137545 0 0 $X=128240 $Y=137355
X48 7 VIA1_C_CDNS_723534627842 $T=130380 81120 0 0 $X=129980 $Y=80930
X49 8 VIA1_C_CDNS_723534627842 $T=132030 81900 0 0 $X=131630 $Y=81710
X50 6 VIA1_C_CDNS_723534627842 $T=134880 137545 0 0 $X=134480 $Y=137355
X51 7 VIA1_C_CDNS_723534627842 $T=137160 81120 0 0 $X=136760 $Y=80930
X52 8 VIA1_C_CDNS_723534627842 $T=137840 81900 0 0 $X=137440 $Y=81710
X53 6 VIA1_C_CDNS_723534627842 $T=141120 137545 0 0 $X=140720 $Y=137355
X54 7 VIA1_C_CDNS_723534627842 $T=142860 81120 0 0 $X=142460 $Y=80930
X55 8 VIA1_C_CDNS_723534627842 $T=144510 81900 0 0 $X=144110 $Y=81710
X56 6 VIA1_C_CDNS_723534627842 $T=147360 137545 0 0 $X=146960 $Y=137355
X57 7 VIA1_C_CDNS_723534627842 $T=149640 81120 0 0 $X=149240 $Y=80930
X58 8 VIA1_C_CDNS_723534627842 $T=150320 81900 0 0 $X=149920 $Y=81710
X59 6 VIA1_C_CDNS_723534627842 $T=153600 137545 0 0 $X=153200 $Y=137355
X60 7 VIA1_C_CDNS_723534627842 $T=155340 81120 0 0 $X=154940 $Y=80930
X61 8 VIA1_C_CDNS_723534627842 $T=156990 81900 0 0 $X=156590 $Y=81710
X62 6 VIA1_C_CDNS_723534627842 $T=159840 137545 0 0 $X=159440 $Y=137355
X63 7 VIA1_C_CDNS_723534627842 $T=162120 81120 0 0 $X=161720 $Y=80930
X64 8 VIA1_C_CDNS_723534627842 $T=162800 81900 0 0 $X=162400 $Y=81710
X65 6 VIA1_C_CDNS_723534627842 $T=166080 137545 0 0 $X=165680 $Y=137355
X66 7 VIA1_C_CDNS_723534627842 $T=167820 81120 0 0 $X=167420 $Y=80930
X67 8 VIA1_C_CDNS_723534627842 $T=169470 81900 0 0 $X=169070 $Y=81710
X68 6 VIA1_C_CDNS_723534627842 $T=172320 137545 0 0 $X=171920 $Y=137355
X69 7 VIA1_C_CDNS_723534627842 $T=174600 81120 0 0 $X=174200 $Y=80930
X70 8 VIA1_C_CDNS_723534627842 $T=175280 81900 0 0 $X=174880 $Y=81710
X71 6 VIA1_C_CDNS_723534627842 $T=178560 137545 0 0 $X=178160 $Y=137355
X72 7 VIA1_C_CDNS_723534627842 $T=180300 81120 0 0 $X=179900 $Y=80930
X73 8 VIA1_C_CDNS_723534627842 $T=181950 81900 0 0 $X=181550 $Y=81710
X74 6 VIA1_C_CDNS_723534627842 $T=184800 137545 0 0 $X=184400 $Y=137355
X75 7 VIA1_C_CDNS_723534627842 $T=187080 81120 0 0 $X=186680 $Y=80930
X76 8 VIA1_C_CDNS_723534627842 $T=187760 81900 0 0 $X=187360 $Y=81710
X77 6 VIA1_C_CDNS_723534627842 $T=191040 137545 0 0 $X=190640 $Y=137355
X78 7 VIA1_C_CDNS_723534627842 $T=192780 81120 0 0 $X=192380 $Y=80930
X79 8 VIA1_C_CDNS_723534627842 $T=194430 81900 0 0 $X=194030 $Y=81710
X80 6 VIA1_C_CDNS_723534627842 $T=197280 137545 0 0 $X=196880 $Y=137355
X81 7 VIA1_C_CDNS_723534627842 $T=199560 81120 0 0 $X=199160 $Y=80930
X82 8 VIA1_C_CDNS_723534627842 $T=200240 81900 0 0 $X=199840 $Y=81710
X83 11 VIA1_C_CDNS_723534627842 $T=248180 27500 0 0 $X=247780 $Y=27310
X84 11 VIA1_C_CDNS_723534627842 $T=249410 27500 0 0 $X=249010 $Y=27310
X85 11 VIA1_C_CDNS_723534627842 $T=250450 27500 0 0 $X=250050 $Y=27310
X86 11 VIA1_C_CDNS_723534627842 $T=251680 27500 0 0 $X=251280 $Y=27310
X87 1 VIA2_C_CDNS_723534627843 $T=8380 17610 0 0 $X=7410 $Y=16950
X88 1 VIA2_C_CDNS_723534627843 $T=8380 49670 0 0 $X=7410 $Y=49010
X89 3 VIA2_C_CDNS_723534627843 $T=10660 15770 0 0 $X=9690 $Y=15110
X90 3 VIA2_C_CDNS_723534627843 $T=10660 47830 0 0 $X=9690 $Y=47170
X91 5 VIA2_C_CDNS_723534627843 $T=12940 13930 0 0 $X=11970 $Y=13270
X92 5 VIA2_C_CDNS_723534627843 $T=12940 45990 0 0 $X=11970 $Y=45330
X93 3 VIA2_C_CDNS_723534627843 $T=76860 15770 0 0 $X=75890 $Y=15110
X94 3 VIA2_C_CDNS_723534627843 $T=76860 47830 0 0 $X=75890 $Y=47170
X95 5 VIA2_C_CDNS_723534627843 $T=79200 13930 0 0 $X=78230 $Y=13270
X96 5 VIA2_C_CDNS_723534627843 $T=79200 45990 0 0 $X=78230 $Y=45330
X97 1 VIA2_C_CDNS_723534627843 $T=81540 17610 0 0 $X=80570 $Y=16950
X98 1 VIA2_C_CDNS_723534627843 $T=81540 49670 0 0 $X=80570 $Y=49010
X99 11 VIA2_C_CDNS_723534627843 $T=102350 65860 0 0 $X=101380 $Y=65200
X100 11 VIA2_C_CDNS_723534627843 $T=102350 98940 0 0 $X=101380 $Y=98280
X101 6 VIA2_C_CDNS_723534627843 $T=104030 116805 0 0 $X=103060 $Y=116145
X102 6 VIA2_C_CDNS_723534627843 $T=104030 158145 0 0 $X=103060 $Y=157485
X103 12 VIA2_C_CDNS_723534627843 $T=104630 64080 0 0 $X=103660 $Y=63420
X104 12 VIA2_C_CDNS_723534627843 $T=104630 97160 0 0 $X=103660 $Y=96500
X105 7 VIA2_C_CDNS_723534627843 $T=106310 120365 0 0 $X=105340 $Y=119705
X106 7 VIA2_C_CDNS_723534627843 $T=106310 152805 0 0 $X=105340 $Y=152145
X107 13 VIA2_C_CDNS_723534627843 $T=106910 67640 0 0 $X=105940 $Y=66980
X108 13 VIA2_C_CDNS_723534627843 $T=106910 95380 0 0 $X=105940 $Y=94720
X109 13 VIA2_C_CDNS_723534627843 $T=108590 118585 0 0 $X=107620 $Y=117925
X110 13 VIA2_C_CDNS_723534627843 $T=108590 156365 0 0 $X=107620 $Y=155705
X111 14 VIA2_C_CDNS_723534627843 $T=110870 123925 0 0 $X=109900 $Y=123265
X112 14 VIA2_C_CDNS_723534627843 $T=110870 151025 0 0 $X=109900 $Y=150365
X113 14 VIA2_C_CDNS_723534627843 $T=208810 123925 0 0 $X=207840 $Y=123265
X114 14 VIA2_C_CDNS_723534627843 $T=208810 151025 0 0 $X=207840 $Y=150365
X115 13 VIA2_C_CDNS_723534627843 $T=211090 67640 0 0 $X=210120 $Y=66980
X116 13 VIA2_C_CDNS_723534627843 $T=211090 95380 0 0 $X=210120 $Y=94720
X117 13 VIA2_C_CDNS_723534627843 $T=211090 118585 0 0 $X=210120 $Y=117925
X118 13 VIA2_C_CDNS_723534627843 $T=211090 156365 0 0 $X=210120 $Y=155705
X119 11 VIA2_C_CDNS_723534627843 $T=213370 65860 0 0 $X=212400 $Y=65200
X120 11 VIA2_C_CDNS_723534627843 $T=213370 98940 0 0 $X=212400 $Y=98280
X121 8 VIA2_C_CDNS_723534627843 $T=213370 122145 0 0 $X=212400 $Y=121485
X122 8 VIA2_C_CDNS_723534627843 $T=213370 154585 0 0 $X=212400 $Y=153925
X123 12 VIA2_C_CDNS_723534627843 $T=215650 64080 0 0 $X=214680 $Y=63420
X124 12 VIA2_C_CDNS_723534627843 $T=215650 97160 0 0 $X=214680 $Y=96500
X125 6 VIA2_C_CDNS_723534627843 $T=215650 116805 0 0 $X=214680 $Y=116145
X126 6 VIA2_C_CDNS_723534627843 $T=215650 158145 0 0 $X=214680 $Y=157485
X127 11 VIA2_C_CDNS_723534627843 $T=227815 16050 0 0 $X=226845 $Y=15390
X128 11 VIA2_C_CDNS_723534627843 $T=227815 37420 0 0 $X=226845 $Y=36760
X129 12 VIA2_C_CDNS_723534627843 $T=239775 17830 0 0 $X=238805 $Y=17170
X130 12 VIA2_C_CDNS_723534627843 $T=239775 35640 0 0 $X=238805 $Y=34980
X131 3 VIA2_C_CDNS_723534627844 $T=44040 62810 0 0 $X=41990 $Y=62060
X132 5 VIA2_C_CDNS_723534627844 $T=78860 62950 0 0 $X=76810 $Y=62200
X133 15 VIA2_C_CDNS_723534627844 $T=311195 26360 0 0 $X=309145 $Y=25610
X134 16 VIA2_C_CDNS_723534627844 $T=315635 26360 0 0 $X=313585 $Y=25610
X135 15 VIA2_C_CDNS_723534627844 $T=324920 82035 0 0 $X=322870 $Y=81285
X136 1 VIA2_C_CDNS_723534627845 $T=8380 31900 0 0 $X=7410 $Y=31760
X137 1 VIA2_C_CDNS_723534627845 $T=81540 31900 0 0 $X=80570 $Y=31760
X138 6 VIA2_C_CDNS_723534627845 $T=104030 137545 0 0 $X=103060 $Y=137405
X139 6 VIA2_C_CDNS_723534627845 $T=215650 137545 0 0 $X=214680 $Y=137405
X140 9 VIA1_C_CDNS_723534627846 $T=15280 19450 0 0 $X=14310 $Y=18790
X141 9 VIA1_C_CDNS_723534627846 $T=15280 44150 0 0 $X=14310 $Y=43490
X142 9 VIA1_C_CDNS_723534627846 $T=74520 19450 0 0 $X=73550 $Y=18790
X143 9 VIA1_C_CDNS_723534627846 $T=74520 44150 0 0 $X=73550 $Y=43490
X144 9 VIA1_C_CDNS_723534627846 $T=230095 19610 0 0 $X=229125 $Y=18950
X145 9 VIA1_C_CDNS_723534627846 $T=230095 33860 0 0 $X=229125 $Y=33200
X146 9 VIA1_C_CDNS_723534627846 $T=237495 19610 0 0 $X=236525 $Y=18950
X147 9 VIA1_C_CDNS_723534627846 $T=237495 33860 0 0 $X=236525 $Y=33200
X148 12 VIA1_C_CDNS_723534627847 $T=201995 64080 0 0 $X=201545 $Y=63680
X149 11 VIA1_C_CDNS_723534627847 $T=201995 98940 0 0 $X=201545 $Y=98540
X150 13 VIA1_C_CDNS_723534627848 $T=115670 67640 0 0 $X=115480 $Y=66980
X151 13 VIA1_C_CDNS_723534627848 $T=115670 95380 0 0 $X=115480 $Y=94720
X152 11 VIA1_C_CDNS_723534627848 $T=121210 65860 0 0 $X=121020 $Y=65200
X153 12 VIA1_C_CDNS_723534627848 $T=121210 97160 0 0 $X=121020 $Y=96500
X154 13 VIA1_C_CDNS_723534627848 $T=121910 67640 0 0 $X=121720 $Y=66980
X155 13 VIA1_C_CDNS_723534627848 $T=121910 95380 0 0 $X=121720 $Y=94720
X156 12 VIA1_C_CDNS_723534627848 $T=127450 64080 0 0 $X=127260 $Y=63420
X157 11 VIA1_C_CDNS_723534627848 $T=127450 98940 0 0 $X=127260 $Y=98280
X158 13 VIA1_C_CDNS_723534627848 $T=128150 67640 0 0 $X=127960 $Y=66980
X159 13 VIA1_C_CDNS_723534627848 $T=128150 95380 0 0 $X=127960 $Y=94720
X160 11 VIA1_C_CDNS_723534627848 $T=133690 65860 0 0 $X=133500 $Y=65200
X161 12 VIA1_C_CDNS_723534627848 $T=133690 97160 0 0 $X=133500 $Y=96500
X162 13 VIA1_C_CDNS_723534627848 $T=134390 67640 0 0 $X=134200 $Y=66980
X163 13 VIA1_C_CDNS_723534627848 $T=134390 95380 0 0 $X=134200 $Y=94720
X164 12 VIA1_C_CDNS_723534627848 $T=139930 64080 0 0 $X=139740 $Y=63420
X165 11 VIA1_C_CDNS_723534627848 $T=139930 98940 0 0 $X=139740 $Y=98280
X166 13 VIA1_C_CDNS_723534627848 $T=140630 67640 0 0 $X=140440 $Y=66980
X167 13 VIA1_C_CDNS_723534627848 $T=140630 95380 0 0 $X=140440 $Y=94720
X168 11 VIA1_C_CDNS_723534627848 $T=146170 65860 0 0 $X=145980 $Y=65200
X169 12 VIA1_C_CDNS_723534627848 $T=146170 97160 0 0 $X=145980 $Y=96500
X170 13 VIA1_C_CDNS_723534627848 $T=146870 67640 0 0 $X=146680 $Y=66980
X171 13 VIA1_C_CDNS_723534627848 $T=146870 95380 0 0 $X=146680 $Y=94720
X172 12 VIA1_C_CDNS_723534627848 $T=152410 64080 0 0 $X=152220 $Y=63420
X173 11 VIA1_C_CDNS_723534627848 $T=152410 98940 0 0 $X=152220 $Y=98280
X174 13 VIA1_C_CDNS_723534627848 $T=153110 67640 0 0 $X=152920 $Y=66980
X175 13 VIA1_C_CDNS_723534627848 $T=153110 95380 0 0 $X=152920 $Y=94720
X176 11 VIA1_C_CDNS_723534627848 $T=158650 65860 0 0 $X=158460 $Y=65200
X177 12 VIA1_C_CDNS_723534627848 $T=158650 97160 0 0 $X=158460 $Y=96500
X178 13 VIA1_C_CDNS_723534627848 $T=159350 67640 0 0 $X=159160 $Y=66980
X179 13 VIA1_C_CDNS_723534627848 $T=159350 95380 0 0 $X=159160 $Y=94720
X180 12 VIA1_C_CDNS_723534627848 $T=164890 64080 0 0 $X=164700 $Y=63420
X181 11 VIA1_C_CDNS_723534627848 $T=164890 98940 0 0 $X=164700 $Y=98280
X182 13 VIA1_C_CDNS_723534627848 $T=165590 67640 0 0 $X=165400 $Y=66980
X183 13 VIA1_C_CDNS_723534627848 $T=165590 95380 0 0 $X=165400 $Y=94720
X184 11 VIA1_C_CDNS_723534627848 $T=171130 65860 0 0 $X=170940 $Y=65200
X185 12 VIA1_C_CDNS_723534627848 $T=171130 97160 0 0 $X=170940 $Y=96500
X186 13 VIA1_C_CDNS_723534627848 $T=171830 67640 0 0 $X=171640 $Y=66980
X187 13 VIA1_C_CDNS_723534627848 $T=171830 95380 0 0 $X=171640 $Y=94720
X188 12 VIA1_C_CDNS_723534627848 $T=177370 64080 0 0 $X=177180 $Y=63420
X189 11 VIA1_C_CDNS_723534627848 $T=177370 98940 0 0 $X=177180 $Y=98280
X190 13 VIA1_C_CDNS_723534627848 $T=178070 67640 0 0 $X=177880 $Y=66980
X191 13 VIA1_C_CDNS_723534627848 $T=178070 95380 0 0 $X=177880 $Y=94720
X192 11 VIA1_C_CDNS_723534627848 $T=183610 65860 0 0 $X=183420 $Y=65200
X193 12 VIA1_C_CDNS_723534627848 $T=183610 97160 0 0 $X=183420 $Y=96500
X194 13 VIA1_C_CDNS_723534627848 $T=184310 67640 0 0 $X=184120 $Y=66980
X195 13 VIA1_C_CDNS_723534627848 $T=184310 95380 0 0 $X=184120 $Y=94720
X196 12 VIA1_C_CDNS_723534627848 $T=189850 64080 0 0 $X=189660 $Y=63420
X197 11 VIA1_C_CDNS_723534627848 $T=189850 98940 0 0 $X=189660 $Y=98280
X198 13 VIA1_C_CDNS_723534627848 $T=190550 67640 0 0 $X=190360 $Y=66980
X199 13 VIA1_C_CDNS_723534627848 $T=190550 95380 0 0 $X=190360 $Y=94720
X200 11 VIA1_C_CDNS_723534627848 $T=196090 65860 0 0 $X=195900 $Y=65200
X201 12 VIA1_C_CDNS_723534627848 $T=196090 97160 0 0 $X=195900 $Y=96500
X202 13 VIA1_C_CDNS_723534627848 $T=196790 67640 0 0 $X=196600 $Y=66980
X203 13 VIA1_C_CDNS_723534627848 $T=196790 95380 0 0 $X=196600 $Y=94720
X204 9 VIA1_C_CDNS_723534627849 $T=17150 19450 0 0 $X=17010 $Y=18740
X205 9 VIA1_C_CDNS_723534627849 $T=17150 44150 0 0 $X=17010 $Y=43440
X206 9 VIA1_C_CDNS_723534627849 $T=27690 19450 0 0 $X=27550 $Y=18740
X207 9 VIA1_C_CDNS_723534627849 $T=27690 44150 0 0 $X=27550 $Y=43440
X208 9 VIA1_C_CDNS_723534627849 $T=28390 19450 0 0 $X=28250 $Y=18740
X209 9 VIA1_C_CDNS_723534627849 $T=28390 44150 0 0 $X=28250 $Y=43440
X210 5 VIA1_C_CDNS_723534627849 $T=38930 13930 0 0 $X=38790 $Y=13220
X211 5 VIA1_C_CDNS_723534627849 $T=38930 45990 0 0 $X=38790 $Y=45280
X212 9 VIA1_C_CDNS_723534627849 $T=39630 19450 0 0 $X=39490 $Y=18740
X213 9 VIA1_C_CDNS_723534627849 $T=39630 44150 0 0 $X=39490 $Y=43440
X214 1 VIA1_C_CDNS_723534627849 $T=50170 17610 0 0 $X=50030 $Y=16900
X215 1 VIA1_C_CDNS_723534627849 $T=50170 49670 0 0 $X=50030 $Y=48960
X216 9 VIA1_C_CDNS_723534627849 $T=50870 19450 0 0 $X=50730 $Y=18740
X217 9 VIA1_C_CDNS_723534627849 $T=50870 44150 0 0 $X=50730 $Y=43440
X218 3 VIA1_C_CDNS_723534627849 $T=61410 15770 0 0 $X=61270 $Y=15060
X219 3 VIA1_C_CDNS_723534627849 $T=61410 47830 0 0 $X=61270 $Y=47120
X220 9 VIA1_C_CDNS_723534627849 $T=62110 19450 0 0 $X=61970 $Y=18740
X221 9 VIA1_C_CDNS_723534627849 $T=62110 44150 0 0 $X=61970 $Y=43440
X222 10 VIA1_C_CDNS_723534627849 $T=62695 100410 0 0 $X=62555 $Y=99700
X223 14 VIA1_C_CDNS_723534627849 $T=64235 96850 0 0 $X=64095 $Y=96140
X224 10 VIA1_C_CDNS_723534627849 $T=64935 100410 0 0 $X=64795 $Y=99700
X225 14 VIA1_C_CDNS_723534627849 $T=66475 96850 0 0 $X=66335 $Y=96140
X226 4 VIA1_C_CDNS_723534627849 $T=67175 98630 0 0 $X=67035 $Y=97920
X227 14 VIA1_C_CDNS_723534627849 $T=68715 96850 0 0 $X=68575 $Y=96140
X228 10 VIA1_C_CDNS_723534627849 $T=69415 100410 0 0 $X=69275 $Y=99700
X229 14 VIA1_C_CDNS_723534627849 $T=70955 96850 0 0 $X=70815 $Y=96140
X230 10 VIA1_C_CDNS_723534627849 $T=71655 100410 0 0 $X=71515 $Y=99700
X231 9 VIA1_C_CDNS_723534627849 $T=72650 19450 0 0 $X=72510 $Y=18740
X232 9 VIA1_C_CDNS_723534627849 $T=72650 44150 0 0 $X=72510 $Y=43440
X233 14 VIA1_C_CDNS_723534627849 $T=73195 96850 0 0 $X=73055 $Y=96140
X234 14 VIA1_C_CDNS_723534627849 $T=113390 123925 0 0 $X=113250 $Y=123215
X235 14 VIA1_C_CDNS_723534627849 $T=113390 151025 0 0 $X=113250 $Y=150315
X236 14 VIA1_C_CDNS_723534627849 $T=118930 123925 0 0 $X=118790 $Y=123215
X237 14 VIA1_C_CDNS_723534627849 $T=118930 151025 0 0 $X=118790 $Y=150315
X238 14 VIA1_C_CDNS_723534627849 $T=119630 123925 0 0 $X=119490 $Y=123215
X239 14 VIA1_C_CDNS_723534627849 $T=119630 151025 0 0 $X=119490 $Y=150315
X240 13 VIA1_C_CDNS_723534627849 $T=125170 118585 0 0 $X=125030 $Y=117875
X241 13 VIA1_C_CDNS_723534627849 $T=125170 156365 0 0 $X=125030 $Y=155655
X242 14 VIA1_C_CDNS_723534627849 $T=125870 123925 0 0 $X=125730 $Y=123215
X243 14 VIA1_C_CDNS_723534627849 $T=125870 151025 0 0 $X=125730 $Y=150315
X244 13 VIA1_C_CDNS_723534627849 $T=131410 118585 0 0 $X=131270 $Y=117875
X245 13 VIA1_C_CDNS_723534627849 $T=131410 156365 0 0 $X=131270 $Y=155655
X246 14 VIA1_C_CDNS_723534627849 $T=132110 123925 0 0 $X=131970 $Y=123215
X247 14 VIA1_C_CDNS_723534627849 $T=132110 151025 0 0 $X=131970 $Y=150315
X248 13 VIA1_C_CDNS_723534627849 $T=137650 118585 0 0 $X=137510 $Y=117875
X249 13 VIA1_C_CDNS_723534627849 $T=137650 156365 0 0 $X=137510 $Y=155655
X250 14 VIA1_C_CDNS_723534627849 $T=138350 123925 0 0 $X=138210 $Y=123215
X251 14 VIA1_C_CDNS_723534627849 $T=138350 151025 0 0 $X=138210 $Y=150315
X252 13 VIA1_C_CDNS_723534627849 $T=143890 118585 0 0 $X=143750 $Y=117875
X253 13 VIA1_C_CDNS_723534627849 $T=143890 156365 0 0 $X=143750 $Y=155655
X254 14 VIA1_C_CDNS_723534627849 $T=144590 123925 0 0 $X=144450 $Y=123215
X255 14 VIA1_C_CDNS_723534627849 $T=144590 151025 0 0 $X=144450 $Y=150315
X256 13 VIA1_C_CDNS_723534627849 $T=150130 118585 0 0 $X=149990 $Y=117875
X257 13 VIA1_C_CDNS_723534627849 $T=150130 156365 0 0 $X=149990 $Y=155655
X258 14 VIA1_C_CDNS_723534627849 $T=150830 123925 0 0 $X=150690 $Y=123215
X259 14 VIA1_C_CDNS_723534627849 $T=150830 151025 0 0 $X=150690 $Y=150315
X260 8 VIA1_C_CDNS_723534627849 $T=156370 122145 0 0 $X=156230 $Y=121435
X261 7 VIA1_C_CDNS_723534627849 $T=156370 152805 0 0 $X=156230 $Y=152095
X262 14 VIA1_C_CDNS_723534627849 $T=157070 123925 0 0 $X=156930 $Y=123215
X263 14 VIA1_C_CDNS_723534627849 $T=157070 151025 0 0 $X=156930 $Y=150315
X264 6 VIA1_C_CDNS_723534627849 $T=162610 116805 0 0 $X=162470 $Y=116095
X265 6 VIA1_C_CDNS_723534627849 $T=162610 158145 0 0 $X=162470 $Y=157435
X266 14 VIA1_C_CDNS_723534627849 $T=163310 123925 0 0 $X=163170 $Y=123215
X267 14 VIA1_C_CDNS_723534627849 $T=163310 151025 0 0 $X=163170 $Y=150315
X268 7 VIA1_C_CDNS_723534627849 $T=168850 120365 0 0 $X=168710 $Y=119655
X269 8 VIA1_C_CDNS_723534627849 $T=168850 154585 0 0 $X=168710 $Y=153875
X270 14 VIA1_C_CDNS_723534627849 $T=169550 123925 0 0 $X=169410 $Y=123215
X271 14 VIA1_C_CDNS_723534627849 $T=169550 151025 0 0 $X=169410 $Y=150315
X272 13 VIA1_C_CDNS_723534627849 $T=175090 118585 0 0 $X=174950 $Y=117875
X273 13 VIA1_C_CDNS_723534627849 $T=175090 156365 0 0 $X=174950 $Y=155655
X274 14 VIA1_C_CDNS_723534627849 $T=175790 123925 0 0 $X=175650 $Y=123215
X275 14 VIA1_C_CDNS_723534627849 $T=175790 151025 0 0 $X=175650 $Y=150315
X276 13 VIA1_C_CDNS_723534627849 $T=181330 118585 0 0 $X=181190 $Y=117875
X277 13 VIA1_C_CDNS_723534627849 $T=181330 156365 0 0 $X=181190 $Y=155655
X278 14 VIA1_C_CDNS_723534627849 $T=182030 123925 0 0 $X=181890 $Y=123215
X279 14 VIA1_C_CDNS_723534627849 $T=182030 151025 0 0 $X=181890 $Y=150315
X280 13 VIA1_C_CDNS_723534627849 $T=187570 118585 0 0 $X=187430 $Y=117875
X281 13 VIA1_C_CDNS_723534627849 $T=187570 156365 0 0 $X=187430 $Y=155655
X282 14 VIA1_C_CDNS_723534627849 $T=188270 123925 0 0 $X=188130 $Y=123215
X283 14 VIA1_C_CDNS_723534627849 $T=188270 151025 0 0 $X=188130 $Y=150315
X284 13 VIA1_C_CDNS_723534627849 $T=193810 118585 0 0 $X=193670 $Y=117875
X285 13 VIA1_C_CDNS_723534627849 $T=193810 156365 0 0 $X=193670 $Y=155655
X286 14 VIA1_C_CDNS_723534627849 $T=194510 123925 0 0 $X=194370 $Y=123215
X287 14 VIA1_C_CDNS_723534627849 $T=194510 151025 0 0 $X=194370 $Y=150315
X288 13 VIA1_C_CDNS_723534627849 $T=200050 118585 0 0 $X=199910 $Y=117875
X289 13 VIA1_C_CDNS_723534627849 $T=200050 156365 0 0 $X=199910 $Y=155655
X290 14 VIA1_C_CDNS_723534627849 $T=200750 123925 0 0 $X=200610 $Y=123215
X291 14 VIA1_C_CDNS_723534627849 $T=200750 151025 0 0 $X=200610 $Y=150315
X292 14 VIA1_C_CDNS_723534627849 $T=206290 123925 0 0 $X=206150 $Y=123215
X293 14 VIA1_C_CDNS_723534627849 $T=206290 151025 0 0 $X=206150 $Y=150315
X294 9 VIA1_C_CDNS_723534627849 $T=231905 19610 0 0 $X=231765 $Y=18900
X295 9 VIA1_C_CDNS_723534627849 $T=231905 33860 0 0 $X=231765 $Y=33150
X296 11 VIA1_C_CDNS_723534627849 $T=233445 16050 0 0 $X=233305 $Y=15340
X297 12 VIA1_C_CDNS_723534627849 $T=233445 35640 0 0 $X=233305 $Y=34930
X298 9 VIA1_C_CDNS_723534627849 $T=234145 19610 0 0 $X=234005 $Y=18900
X299 9 VIA1_C_CDNS_723534627849 $T=234145 33860 0 0 $X=234005 $Y=33150
X300 12 VIA1_C_CDNS_723534627849 $T=235685 17830 0 0 $X=235545 $Y=17120
X301 11 VIA1_C_CDNS_723534627849 $T=235685 37420 0 0 $X=235545 $Y=36710
X302 17 VIA1_C_CDNS_7235346278410 $T=109005 31610 0 0 $X=108815 $Y=31420
X303 18 VIA1_C_CDNS_7235346278410 $T=109625 32170 0 0 $X=109435 $Y=31980
X304 17 VIA1_C_CDNS_7235346278410 $T=114545 31610 0 0 $X=114355 $Y=31420
X305 18 VIA1_C_CDNS_7235346278410 $T=115165 32170 0 0 $X=114975 $Y=31980
X306 17 VIA1_C_CDNS_7235346278410 $T=120085 31610 0 0 $X=119895 $Y=31420
X307 18 VIA1_C_CDNS_7235346278410 $T=120705 32170 0 0 $X=120515 $Y=31980
X308 17 VIA1_C_CDNS_7235346278410 $T=125625 31610 0 0 $X=125435 $Y=31420
X309 18 VIA1_C_CDNS_7235346278410 $T=126245 32170 0 0 $X=126055 $Y=31980
X310 17 VIA1_C_CDNS_7235346278410 $T=131165 31610 0 0 $X=130975 $Y=31420
X311 18 VIA1_C_CDNS_7235346278410 $T=131785 32170 0 0 $X=131595 $Y=31980
X312 17 VIA1_C_CDNS_7235346278410 $T=136705 31610 0 0 $X=136515 $Y=31420
X313 18 VIA1_C_CDNS_7235346278410 $T=137325 32170 0 0 $X=137135 $Y=31980
X314 17 VIA1_C_CDNS_7235346278410 $T=142245 31610 0 0 $X=142055 $Y=31420
X315 18 VIA1_C_CDNS_7235346278410 $T=142865 32170 0 0 $X=142675 $Y=31980
X316 17 VIA1_C_CDNS_7235346278410 $T=147785 31610 0 0 $X=147595 $Y=31420
X317 18 VIA1_C_CDNS_7235346278410 $T=148405 32170 0 0 $X=148215 $Y=31980
X318 17 VIA1_C_CDNS_7235346278410 $T=153325 31610 0 0 $X=153135 $Y=31420
X319 18 VIA1_C_CDNS_7235346278410 $T=153945 32170 0 0 $X=153755 $Y=31980
X320 17 VIA1_C_CDNS_7235346278410 $T=163595 31610 0 0 $X=163405 $Y=31420
X321 18 VIA1_C_CDNS_7235346278410 $T=164105 32170 0 0 $X=163915 $Y=31980
X322 17 VIA1_C_CDNS_7235346278410 $T=169135 31610 0 0 $X=168945 $Y=31420
X323 18 VIA1_C_CDNS_7235346278410 $T=169645 32170 0 0 $X=169455 $Y=31980
X324 17 VIA1_C_CDNS_7235346278410 $T=174675 31610 0 0 $X=174485 $Y=31420
X325 18 VIA1_C_CDNS_7235346278410 $T=175185 32170 0 0 $X=174995 $Y=31980
X326 17 VIA1_C_CDNS_7235346278410 $T=180215 31610 0 0 $X=180025 $Y=31420
X327 18 VIA1_C_CDNS_7235346278410 $T=180725 32170 0 0 $X=180535 $Y=31980
X328 17 VIA1_C_CDNS_7235346278410 $T=185755 31610 0 0 $X=185565 $Y=31420
X329 18 VIA1_C_CDNS_7235346278410 $T=186265 32170 0 0 $X=186075 $Y=31980
X330 17 VIA1_C_CDNS_7235346278410 $T=191295 31610 0 0 $X=191105 $Y=31420
X331 18 VIA1_C_CDNS_7235346278410 $T=191805 32170 0 0 $X=191615 $Y=31980
X332 17 VIA1_C_CDNS_7235346278410 $T=196835 31610 0 0 $X=196645 $Y=31420
X333 18 VIA1_C_CDNS_7235346278410 $T=197345 32170 0 0 $X=197155 $Y=31980
X334 17 VIA1_C_CDNS_7235346278410 $T=202375 31610 0 0 $X=202185 $Y=31420
X335 18 VIA1_C_CDNS_7235346278410 $T=202885 32170 0 0 $X=202695 $Y=31980
X336 17 VIA1_C_CDNS_7235346278410 $T=207915 31610 0 0 $X=207725 $Y=31420
X337 18 VIA1_C_CDNS_7235346278410 $T=208425 32170 0 0 $X=208235 $Y=31980
X338 7 9 ND_C_CDNS_7235346278411 $T=131350 17825 0 0 $X=106195 $Y=17420
X339 8 9 ND_C_CDNS_7235346278411 $T=131350 45950 0 0 $X=106195 $Y=45545
X340 8 9 ND_C_CDNS_7235346278411 $T=185880 16050 0 0 $X=160725 $Y=15645
X341 7 9 ND_C_CDNS_7235346278411 $T=185880 47720 0 0 $X=160725 $Y=47315
X342 9 VIA2_C_CDNS_7235346278412 $T=112085 14270 0 0 $X=111685 $Y=13560
X343 9 VIA2_C_CDNS_7235346278412 $T=112085 49510 0 0 $X=111685 $Y=48800
X344 9 VIA2_C_CDNS_7235346278412 $T=123165 14270 0 0 $X=122765 $Y=13560
X345 9 VIA2_C_CDNS_7235346278412 $T=123165 49510 0 0 $X=122765 $Y=48800
X346 9 VIA2_C_CDNS_7235346278412 $T=134245 14270 0 0 $X=133845 $Y=13560
X347 9 VIA2_C_CDNS_7235346278412 $T=134245 49510 0 0 $X=133845 $Y=48800
X348 9 VIA2_C_CDNS_7235346278412 $T=145325 14270 0 0 $X=144925 $Y=13560
X349 9 VIA2_C_CDNS_7235346278412 $T=145325 49510 0 0 $X=144925 $Y=48800
X350 9 VIA2_C_CDNS_7235346278412 $T=156405 14270 0 0 $X=156005 $Y=13560
X351 9 VIA2_C_CDNS_7235346278412 $T=156405 49510 0 0 $X=156005 $Y=48800
X352 9 VIA2_C_CDNS_7235346278412 $T=166365 14270 0 0 $X=165965 $Y=13560
X353 9 VIA2_C_CDNS_7235346278412 $T=166365 49510 0 0 $X=165965 $Y=48800
X354 9 VIA2_C_CDNS_7235346278412 $T=177445 14270 0 0 $X=177045 $Y=13560
X355 9 VIA2_C_CDNS_7235346278412 $T=177445 49510 0 0 $X=177045 $Y=48800
X356 9 VIA2_C_CDNS_7235346278412 $T=188525 14270 0 0 $X=188125 $Y=13560
X357 9 VIA2_C_CDNS_7235346278412 $T=188525 49510 0 0 $X=188125 $Y=48800
X358 9 VIA2_C_CDNS_7235346278412 $T=199605 14270 0 0 $X=199205 $Y=13560
X359 9 VIA2_C_CDNS_7235346278412 $T=199605 49510 0 0 $X=199205 $Y=48800
X360 9 VIA2_C_CDNS_7235346278412 $T=210685 14270 0 0 $X=210285 $Y=13560
X361 9 VIA2_C_CDNS_7235346278412 $T=210685 49510 0 0 $X=210285 $Y=48800
X362 19 VIA1_C_CDNS_7235346278413 $T=13505 83830 1 0 $X=13015 $Y=83600
X363 19 VIA1_C_CDNS_7235346278413 $T=13505 86055 0 0 $X=13015 $Y=85825
X364 20 VIA1_C_CDNS_7235346278413 $T=17705 83830 1 0 $X=17215 $Y=83600
X365 20 VIA1_C_CDNS_7235346278413 $T=17705 86055 0 0 $X=17215 $Y=85825
X366 21 VIA1_C_CDNS_7235346278414 $T=23615 88310 0 0 $X=22865 $Y=88080
X367 22 VIA1_C_CDNS_7235346278414 $T=24350 86955 0 0 $X=23600 $Y=86725
X368 9 VIA1_C_CDNS_7235346278416 $T=105815 12260 0 0 $X=103025 $Y=11060
X369 9 VIA1_C_CDNS_7235346278416 $T=211445 12030 0 0 $X=208655 $Y=10830
X370 9 VIA2_C_CDNS_7235346278417 $T=105815 12260 0 0 $X=103025 $Y=11060
X371 9 VIA2_C_CDNS_7235346278417 $T=211445 12030 0 0 $X=208655 $Y=10830
X372 7 VIA1_C_CDNS_7235346278418 $T=101790 44390 0 0 $X=101040 $Y=42080
X373 8 VIA1_C_CDNS_7235346278418 $T=215715 44390 0 0 $X=214965 $Y=42080
X374 9 VIA1_C_CDNS_7235346278419 $T=243980 19610 0 0 $X=241930 $Y=18860
X375 15 VIA1_C_CDNS_7235346278419 $T=311195 26360 0 0 $X=309145 $Y=25610
X376 16 VIA1_C_CDNS_7235346278419 $T=315635 26360 0 0 $X=313585 $Y=25610
X377 15 VIA1_C_CDNS_7235346278419 $T=324920 82035 0 0 $X=322870 $Y=81285
X378 10 VIA2_C_CDNS_7235346278420 $T=92185 100410 0 0 $X=89615 $Y=99660
X379 10 VIA2_C_CDNS_7235346278420 $T=249890 17585 0 0 $X=247320 $Y=16835
X380 14 9 VIA2_C_CDNS_7235346278422 $T=110885 161700 0 0 $X=108315 $Y=160170
X381 14 9 VIA2_C_CDNS_7235346278422 $T=208825 161700 0 0 $X=206255 $Y=160170
X382 14 9 VIA1_C_CDNS_7235346278423 $T=105735 160860 0 0 $X=97965 $Y=160110
X383 14 9 VIA1_C_CDNS_7235346278423 $T=213285 160860 0 0 $X=205515 $Y=160110
X384 15 VIA3_C_CDNS_7235346278432 $T=311195 26360 0 0 $X=309145 $Y=25610
X385 16 VIA3_C_CDNS_7235346278432 $T=315635 26360 0 0 $X=313585 $Y=25610
X386 15 VIA3_C_CDNS_7235346278432 $T=324920 82035 0 0 $X=322870 $Y=81285
X387 18 VIA2_C_CDNS_7235346278438 $T=98240 32160 0 0 $X=97490 $Y=31410
X388 10 VIA2_C_CDNS_7235346278438 $T=259885 73765 0 0 $X=259135 $Y=73015
X389 23 VIATP_C_CDNS_7235346278440 $T=376900 51365 0 0 $X=376110 $Y=50835
X390 23 VIATP_C_CDNS_7235346278440 $T=376900 147425 0 0 $X=376110 $Y=146895
X391 24 VIATP_C_CDNS_7235346278440 $T=557055 51365 0 0 $X=556265 $Y=50835
X392 24 VIATP_C_CDNS_7235346278440 $T=557055 147425 0 0 $X=556265 $Y=146895
X393 23 VIATP_C_CDNS_7235346278444 $T=433355 51365 0 0 $X=432695 $Y=50835
X394 23 VIATP_C_CDNS_7235346278444 $T=433355 147425 0 0 $X=432695 $Y=146895
X395 24 VIATP_C_CDNS_7235346278444 $T=500600 51365 0 0 $X=499940 $Y=50835
X396 24 VIATP_C_CDNS_7235346278444 $T=500600 147425 0 0 $X=499940 $Y=146895
X397 19 VIA2_C_CDNS_7235346278453 $T=13245 83830 0 0 $X=12495 $Y=83600
X398 20 VIA2_C_CDNS_7235346278453 $T=17445 83830 0 0 $X=16695 $Y=83600
X399 9 11 10 ne3_CDNS_723534627840 $T=248120 21400 0 0 $X=247320 $Y=21000
X400 25 15 16 10 nedia_CDNS_723534627841 $T=282450 37820 0 0 $X=266230 $Y=18430
X401 9 22 1 ne3_CDNS_723534627842 $T=25060 81535 0 0 $X=24260 $Y=80955
X402 9 21 11 ne3_CDNS_723534627842 $T=30635 81535 0 0 $X=29835 $Y=80955
X403 15 16 25 rpp1k1_3_CDNS_723534627843 $T=317545 27490 0 90 $X=309065 $Y=26550
X404 25 24 23 15 nedia_CDNS_723534627844 $T=441980 141045 0 270 $X=422590 $Y=41525
X405 1 2 2 9 ne3_CDNS_723534627845 $T=8060 64240 0 0 $X=7260 $Y=63840
X406 3 2 4 9 ne3_CDNS_723534627845 $T=33845 64240 0 0 $X=33045 $Y=63840
X407 5 2 6 9 ne3_CDNS_723534627845 $T=59570 64240 0 0 $X=58770 $Y=63840
X408 14 4 10 9 pe3_CDNS_723534627846 $T=63965 94930 0 180 $X=61455 $Y=83900
X409 14 4 10 9 pe3_CDNS_723534627846 $T=66205 94930 0 180 $X=63695 $Y=83900
X410 14 4 4 9 pe3_CDNS_723534627846 $T=68445 94930 0 180 $X=65935 $Y=83900
X411 14 4 10 9 pe3_CDNS_723534627846 $T=70685 94930 0 180 $X=68175 $Y=83900
X412 14 4 10 9 pe3_CDNS_723534627846 $T=72925 94930 0 180 $X=70415 $Y=83900
X413 14 19 22 9 pe3_CDNS_723534627847 $T=15530 89865 0 180 $X=13480 $Y=86295
X414 14 20 21 9 pe3_CDNS_723534627847 $T=19690 89865 0 180 $X=17640 $Y=86295
X415 16 24 25 rpp1k1_3_CDNS_723534627848 $T=558265 45130 0 90 $X=515365 $Y=41970
X416 14 14 14 14 9 pe3_CDNS_7235346278411 $T=109700 69700 0 0 $X=108190 $Y=68670
X417 14 14 14 14 9 pe3_CDNS_7235346278411 $T=109700 93320 1 0 $X=108190 $Y=82290
X418 14 14 14 14 9 pe3_CDNS_7235346278411 $T=113660 125985 0 0 $X=112150 $Y=124955
X419 14 14 14 14 9 pe3_CDNS_7235346278411 $T=113660 148965 1 0 $X=112150 $Y=137935
X420 13 8 11 14 9 pe3_CDNS_7235346278411 $T=115940 69700 0 0 $X=114430 $Y=68670
X421 13 7 12 14 9 pe3_CDNS_7235346278411 $T=115940 93320 1 0 $X=114430 $Y=82290
X422 14 6 13 14 9 pe3_CDNS_7235346278411 $T=119900 125985 0 0 $X=118390 $Y=124955
X423 14 6 13 14 9 pe3_CDNS_7235346278411 $T=119900 148965 1 0 $X=118390 $Y=137935
X424 13 7 12 14 9 pe3_CDNS_7235346278411 $T=122180 69700 0 0 $X=120670 $Y=68670
X425 13 8 11 14 9 pe3_CDNS_7235346278411 $T=122180 93320 1 0 $X=120670 $Y=82290
X426 14 6 13 14 9 pe3_CDNS_7235346278411 $T=126140 125985 0 0 $X=124630 $Y=124955
X427 14 6 13 14 9 pe3_CDNS_7235346278411 $T=126140 148965 1 0 $X=124630 $Y=137935
X428 13 8 11 14 9 pe3_CDNS_7235346278411 $T=128420 69700 0 0 $X=126910 $Y=68670
X429 13 7 12 14 9 pe3_CDNS_7235346278411 $T=128420 93320 1 0 $X=126910 $Y=82290
X430 14 6 13 14 9 pe3_CDNS_7235346278411 $T=132380 125985 0 0 $X=130870 $Y=124955
X431 14 6 13 14 9 pe3_CDNS_7235346278411 $T=132380 148965 1 0 $X=130870 $Y=137935
X432 13 7 12 14 9 pe3_CDNS_7235346278411 $T=134660 69700 0 0 $X=133150 $Y=68670
X433 13 8 11 14 9 pe3_CDNS_7235346278411 $T=134660 93320 1 0 $X=133150 $Y=82290
X434 14 6 13 14 9 pe3_CDNS_7235346278411 $T=138620 125985 0 0 $X=137110 $Y=124955
X435 14 6 13 14 9 pe3_CDNS_7235346278411 $T=138620 148965 1 0 $X=137110 $Y=137935
X436 13 8 11 14 9 pe3_CDNS_7235346278411 $T=140900 69700 0 0 $X=139390 $Y=68670
X437 13 7 12 14 9 pe3_CDNS_7235346278411 $T=140900 93320 1 0 $X=139390 $Y=82290
X438 14 6 13 14 9 pe3_CDNS_7235346278411 $T=144860 125985 0 0 $X=143350 $Y=124955
X439 14 6 13 14 9 pe3_CDNS_7235346278411 $T=144860 148965 1 0 $X=143350 $Y=137935
X440 13 7 12 14 9 pe3_CDNS_7235346278411 $T=147140 69700 0 0 $X=145630 $Y=68670
X441 13 8 11 14 9 pe3_CDNS_7235346278411 $T=147140 93320 1 0 $X=145630 $Y=82290
X442 14 6 8 14 9 pe3_CDNS_7235346278411 $T=151100 125985 0 0 $X=149590 $Y=124955
X443 14 6 7 14 9 pe3_CDNS_7235346278411 $T=151100 148965 1 0 $X=149590 $Y=137935
X444 13 8 11 14 9 pe3_CDNS_7235346278411 $T=153380 69700 0 0 $X=151870 $Y=68670
X445 13 7 12 14 9 pe3_CDNS_7235346278411 $T=153380 93320 1 0 $X=151870 $Y=82290
X446 14 6 6 14 9 pe3_CDNS_7235346278411 $T=157340 125985 0 0 $X=155830 $Y=124955
X447 14 6 6 14 9 pe3_CDNS_7235346278411 $T=157340 148965 1 0 $X=155830 $Y=137935
X448 13 7 12 14 9 pe3_CDNS_7235346278411 $T=159620 69700 0 0 $X=158110 $Y=68670
X449 13 8 11 14 9 pe3_CDNS_7235346278411 $T=159620 93320 1 0 $X=158110 $Y=82290
X450 14 6 7 14 9 pe3_CDNS_7235346278411 $T=163580 125985 0 0 $X=162070 $Y=124955
X451 14 6 8 14 9 pe3_CDNS_7235346278411 $T=163580 148965 1 0 $X=162070 $Y=137935
X452 13 8 11 14 9 pe3_CDNS_7235346278411 $T=165860 69700 0 0 $X=164350 $Y=68670
X453 13 7 12 14 9 pe3_CDNS_7235346278411 $T=165860 93320 1 0 $X=164350 $Y=82290
X454 14 6 13 14 9 pe3_CDNS_7235346278411 $T=169820 125985 0 0 $X=168310 $Y=124955
X455 14 6 13 14 9 pe3_CDNS_7235346278411 $T=169820 148965 1 0 $X=168310 $Y=137935
X456 13 7 12 14 9 pe3_CDNS_7235346278411 $T=172100 69700 0 0 $X=170590 $Y=68670
X457 13 8 11 14 9 pe3_CDNS_7235346278411 $T=172100 93320 1 0 $X=170590 $Y=82290
X458 14 6 13 14 9 pe3_CDNS_7235346278411 $T=176060 125985 0 0 $X=174550 $Y=124955
X459 14 6 13 14 9 pe3_CDNS_7235346278411 $T=176060 148965 1 0 $X=174550 $Y=137935
X460 13 8 11 14 9 pe3_CDNS_7235346278411 $T=178340 69700 0 0 $X=176830 $Y=68670
X461 13 7 12 14 9 pe3_CDNS_7235346278411 $T=178340 93320 1 0 $X=176830 $Y=82290
X462 14 6 13 14 9 pe3_CDNS_7235346278411 $T=182300 125985 0 0 $X=180790 $Y=124955
X463 14 6 13 14 9 pe3_CDNS_7235346278411 $T=182300 148965 1 0 $X=180790 $Y=137935
X464 13 7 12 14 9 pe3_CDNS_7235346278411 $T=184580 69700 0 0 $X=183070 $Y=68670
X465 13 8 11 14 9 pe3_CDNS_7235346278411 $T=184580 93320 1 0 $X=183070 $Y=82290
X466 14 6 13 14 9 pe3_CDNS_7235346278411 $T=188540 125985 0 0 $X=187030 $Y=124955
X467 14 6 13 14 9 pe3_CDNS_7235346278411 $T=188540 148965 1 0 $X=187030 $Y=137935
X468 13 8 11 14 9 pe3_CDNS_7235346278411 $T=190820 69700 0 0 $X=189310 $Y=68670
X469 13 7 12 14 9 pe3_CDNS_7235346278411 $T=190820 93320 1 0 $X=189310 $Y=82290
X470 14 6 13 14 9 pe3_CDNS_7235346278411 $T=194780 125985 0 0 $X=193270 $Y=124955
X471 14 6 13 14 9 pe3_CDNS_7235346278411 $T=194780 148965 1 0 $X=193270 $Y=137935
X472 13 7 12 14 9 pe3_CDNS_7235346278411 $T=197060 69700 0 0 $X=195550 $Y=68670
X473 13 8 11 14 9 pe3_CDNS_7235346278411 $T=197060 93320 1 0 $X=195550 $Y=82290
X474 14 14 14 14 9 pe3_CDNS_7235346278411 $T=201020 125985 0 0 $X=199510 $Y=124955
X475 14 14 14 14 9 pe3_CDNS_7235346278411 $T=201020 148965 1 0 $X=199510 $Y=137935
X476 14 14 14 14 9 pe3_CDNS_7235346278411 $T=203300 69700 0 0 $X=201790 $Y=68670
X477 14 14 14 14 9 pe3_CDNS_7235346278411 $T=203300 93320 1 0 $X=201790 $Y=82290
X478 9 9 9 ne3_CDNS_7235346278412 $T=17420 20740 0 0 $X=16620 $Y=20340
X479 9 9 9 ne3_CDNS_7235346278412 $T=17420 42860 1 0 $X=16620 $Y=32290
X480 9 1 5 ne3_CDNS_7235346278412 $T=28660 20740 0 0 $X=27860 $Y=20340
X481 9 1 5 ne3_CDNS_7235346278412 $T=28660 42860 1 0 $X=27860 $Y=32290
X482 9 1 1 ne3_CDNS_7235346278412 $T=39900 20740 0 0 $X=39100 $Y=20340
X483 9 1 1 ne3_CDNS_7235346278412 $T=39900 42860 1 0 $X=39100 $Y=32290
X484 9 1 3 ne3_CDNS_7235346278412 $T=51140 20740 0 0 $X=50340 $Y=20340
X485 9 1 3 ne3_CDNS_7235346278412 $T=51140 42860 1 0 $X=50340 $Y=32290
X486 9 9 9 ne3_CDNS_7235346278412 $T=62380 20740 0 0 $X=61580 $Y=20340
X487 9 9 9 ne3_CDNS_7235346278412 $T=62380 42860 1 0 $X=61580 $Y=32290
X488 9 12 11 ne3_CDNS_7235346278413 $T=232175 21040 0 0 $X=231375 $Y=20640
X489 9 12 12 ne3_CDNS_7235346278413 $T=232175 32430 1 0 $X=231375 $Y=26860
X490 9 12 12 ne3_CDNS_7235346278413 $T=234415 21040 0 0 $X=233615 $Y=20640
X491 9 12 11 ne3_CDNS_7235346278413 $T=234415 32430 1 0 $X=233615 $Y=26860
X492 7 18 9 pe3_CDNS_7235346278414 $T=106815 19890 0 0 $X=105305 $Y=18860
X493 8 17 9 pe3_CDNS_7235346278414 $T=106815 43890 1 0 $X=105305 $Y=32860
X494 8 17 9 pe3_CDNS_7235346278414 $T=161095 19890 0 0 $X=159585 $Y=18860
X495 7 18 9 pe3_CDNS_7235346278414 $T=161095 43890 1 0 $X=159585 $Y=32860
X496 23 17 9 rpp1k1_3_CDNS_7235346278415 $T=229190 61300 0 90 $X=226970 $Y=60360
X497 23 17 9 rpp1k1_3_CDNS_7235346278415 $T=232060 61300 0 90 $X=229840 $Y=60360
X498 23 17 9 rpp1k1_3_CDNS_7235346278415 $T=234930 61300 0 90 $X=232710 $Y=60360
X499 23 17 9 rpp1k1_3_CDNS_7235346278415 $T=237800 61300 0 90 $X=235580 $Y=60360
X500 23 17 9 rpp1k1_3_CDNS_7235346278415 $T=240670 61300 0 90 $X=238450 $Y=60360
X501 23 17 9 rpp1k1_3_CDNS_7235346278415 $T=243540 61300 0 90 $X=241320 $Y=60360
X502 23 17 9 rpp1k1_3_CDNS_7235346278415 $T=246410 61300 0 90 $X=244190 $Y=60360
X503 23 17 9 rpp1k1_3_CDNS_7235346278415 $T=249280 61300 0 90 $X=247060 $Y=60360
X504 23 17 9 rpp1k1_3_CDNS_7235346278415 $T=252150 61300 0 90 $X=249930 $Y=60360
X505 10 26 14 9 rpp1k1_3_CDNS_7235346278416 $T=255085 124550 0 180 $X=228430 $Y=99030
X506 27 15 25 rpp1k1_3_CDNS_7235346278417 $T=322885 76685 0 270 $X=322665 $Y=25845
X507 9 19 22 ne3_CDNS_7235346278418 $T=14340 81020 0 0 $X=13540 $Y=80620
X508 9 20 21 ne3_CDNS_7235346278418 $T=18500 81020 0 0 $X=17700 $Y=80620
X509 23 MASCO__X1 $T=432695 51895 0 0 $X=432695 $Y=51895
X510 23 MASCO__X1 $T=432695 56895 0 0 $X=432695 $Y=56895
X511 23 MASCO__X1 $T=432695 61895 0 0 $X=432695 $Y=61895
X512 23 MASCO__X1 $T=432695 66895 0 0 $X=432695 $Y=66895
X513 23 MASCO__X1 $T=432695 71895 0 0 $X=432695 $Y=71895
X514 23 MASCO__X1 $T=432695 76895 0 0 $X=432695 $Y=76895
X515 23 MASCO__X1 $T=432695 81895 0 0 $X=432695 $Y=81895
X516 23 MASCO__X1 $T=432695 86895 0 0 $X=432695 $Y=86895
X517 23 MASCO__X1 $T=432695 91895 0 0 $X=432695 $Y=91895
X518 23 MASCO__X1 $T=432695 96895 0 0 $X=432695 $Y=96895
X519 23 MASCO__X1 $T=432695 101895 0 0 $X=432695 $Y=101895
X520 23 MASCO__X1 $T=432695 106895 0 0 $X=432695 $Y=106895
X521 23 MASCO__X1 $T=432695 111895 0 0 $X=432695 $Y=111895
X522 23 MASCO__X1 $T=432695 116895 0 0 $X=432695 $Y=116895
X523 23 MASCO__X1 $T=432695 121895 0 0 $X=432695 $Y=121895
X524 23 MASCO__X1 $T=432695 126895 0 0 $X=432695 $Y=126895
X525 23 MASCO__X1 $T=432695 131895 0 0 $X=432695 $Y=131895
X526 23 MASCO__X1 $T=432695 136895 0 0 $X=432695 $Y=136895
X527 23 MASCO__X1 $T=432695 141895 0 0 $X=432695 $Y=141895
X528 24 MASCO__X1 $T=499940 51895 0 0 $X=499940 $Y=51895
X529 24 MASCO__X1 $T=499940 56895 0 0 $X=499940 $Y=56895
X530 24 MASCO__X1 $T=499940 61895 0 0 $X=499940 $Y=61895
X531 24 MASCO__X1 $T=499940 66895 0 0 $X=499940 $Y=66895
X532 24 MASCO__X1 $T=499940 71895 0 0 $X=499940 $Y=71895
X533 24 MASCO__X1 $T=499940 76895 0 0 $X=499940 $Y=76895
X534 24 MASCO__X1 $T=499940 81895 0 0 $X=499940 $Y=81895
X535 24 MASCO__X1 $T=499940 86895 0 0 $X=499940 $Y=86895
X536 24 MASCO__X1 $T=499940 91895 0 0 $X=499940 $Y=91895
X537 24 MASCO__X1 $T=499940 96895 0 0 $X=499940 $Y=96895
X538 24 MASCO__X1 $T=499940 101895 0 0 $X=499940 $Y=101895
X539 24 MASCO__X1 $T=499940 106895 0 0 $X=499940 $Y=106895
X540 24 MASCO__X1 $T=499940 111895 0 0 $X=499940 $Y=111895
X541 24 MASCO__X1 $T=499940 116895 0 0 $X=499940 $Y=116895
X542 24 MASCO__X1 $T=499940 121895 0 0 $X=499940 $Y=121895
X543 24 MASCO__X1 $T=499940 126895 0 0 $X=499940 $Y=126895
X544 24 MASCO__X1 $T=499940 131895 0 0 $X=499940 $Y=131895
X545 24 MASCO__X1 $T=499940 136895 0 0 $X=499940 $Y=136895
X546 24 MASCO__X1 $T=499940 141895 0 0 $X=499940 $Y=141895
X547 23 MASCO__X2 $T=376110 51895 0 0 $X=376110 $Y=51895
X548 23 MASCO__X2 $T=376110 56895 0 0 $X=376110 $Y=56895
X549 23 MASCO__X2 $T=376110 61895 0 0 $X=376110 $Y=61895
X550 23 MASCO__X2 $T=376110 66895 0 0 $X=376110 $Y=66895
X551 23 MASCO__X2 $T=376110 71895 0 0 $X=376110 $Y=71895
X552 23 MASCO__X2 $T=376110 76895 0 0 $X=376110 $Y=76895
X553 23 MASCO__X2 $T=376110 81895 0 0 $X=376110 $Y=81895
X554 23 MASCO__X2 $T=376110 86895 0 0 $X=376110 $Y=86895
X555 23 MASCO__X2 $T=376110 91895 0 0 $X=376110 $Y=91895
X556 23 MASCO__X2 $T=376110 96895 0 0 $X=376110 $Y=96895
X557 23 MASCO__X2 $T=376110 101895 0 0 $X=376110 $Y=101895
X558 23 MASCO__X2 $T=376110 106895 0 0 $X=376110 $Y=106895
X559 23 MASCO__X2 $T=376110 111895 0 0 $X=376110 $Y=111895
X560 23 MASCO__X2 $T=376110 116895 0 0 $X=376110 $Y=116895
X561 23 MASCO__X2 $T=376110 121895 0 0 $X=376110 $Y=121895
X562 23 MASCO__X2 $T=376110 126895 0 0 $X=376110 $Y=126895
X563 23 MASCO__X2 $T=376110 131895 0 0 $X=376110 $Y=131895
X564 23 MASCO__X2 $T=376110 136895 0 0 $X=376110 $Y=136895
X565 23 MASCO__X2 $T=376110 141895 0 0 $X=376110 $Y=141895
X566 24 MASCO__X2 $T=556265 51895 0 0 $X=556265 $Y=51895
X567 24 MASCO__X2 $T=556265 56895 0 0 $X=556265 $Y=56895
X568 24 MASCO__X2 $T=556265 61895 0 0 $X=556265 $Y=61895
X569 24 MASCO__X2 $T=556265 66895 0 0 $X=556265 $Y=66895
X570 24 MASCO__X2 $T=556265 71895 0 0 $X=556265 $Y=71895
X571 24 MASCO__X2 $T=556265 76895 0 0 $X=556265 $Y=76895
X572 24 MASCO__X2 $T=556265 81895 0 0 $X=556265 $Y=81895
X573 24 MASCO__X2 $T=556265 86895 0 0 $X=556265 $Y=86895
X574 24 MASCO__X2 $T=556265 91895 0 0 $X=556265 $Y=91895
X575 24 MASCO__X2 $T=556265 96895 0 0 $X=556265 $Y=96895
X576 24 MASCO__X2 $T=556265 101895 0 0 $X=556265 $Y=101895
X577 24 MASCO__X2 $T=556265 106895 0 0 $X=556265 $Y=106895
X578 24 MASCO__X2 $T=556265 111895 0 0 $X=556265 $Y=111895
X579 24 MASCO__X2 $T=556265 116895 0 0 $X=556265 $Y=116895
X580 24 MASCO__X2 $T=556265 121895 0 0 $X=556265 $Y=121895
X581 24 MASCO__X2 $T=556265 126895 0 0 $X=556265 $Y=126895
X582 24 MASCO__X2 $T=556265 131895 0 0 $X=556265 $Y=131895
X583 24 MASCO__X2 $T=556265 136895 0 0 $X=556265 $Y=136895
X584 24 MASCO__X2 $T=556265 141895 0 0 $X=556265 $Y=141895
X585 23 MASCO__Y6 $T=377695 50835 0 0 $X=377695 $Y=50835
X586 23 MASCO__Y6 $T=377695 146895 0 0 $X=377695 $Y=146895
X587 23 MASCO__Y6 $T=388695 50835 0 0 $X=388695 $Y=50835
X588 23 MASCO__Y6 $T=388695 146895 0 0 $X=388695 $Y=146895
X589 23 MASCO__Y6 $T=399695 50835 0 0 $X=399695 $Y=50835
X590 23 MASCO__Y6 $T=399695 146895 0 0 $X=399695 $Y=146895
X591 23 MASCO__Y6 $T=410695 50835 0 0 $X=410695 $Y=50835
X592 23 MASCO__Y6 $T=410695 146895 0 0 $X=410695 $Y=146895
X593 23 MASCO__Y6 $T=421695 50835 0 0 $X=421695 $Y=50835
X594 23 MASCO__Y6 $T=421695 146895 0 0 $X=421695 $Y=146895
X595 24 MASCO__Y6 $T=501265 50835 0 0 $X=501265 $Y=50835
X596 24 MASCO__Y6 $T=501265 146895 0 0 $X=501265 $Y=146895
X597 24 MASCO__Y6 $T=512265 50835 0 0 $X=512265 $Y=50835
X598 24 MASCO__Y6 $T=512265 146895 0 0 $X=512265 $Y=146895
X599 24 MASCO__Y6 $T=523265 50835 0 0 $X=523265 $Y=50835
X600 24 MASCO__Y6 $T=523265 146895 0 0 $X=523265 $Y=146895
X601 24 MASCO__Y6 $T=534265 50835 0 0 $X=534265 $Y=50835
X602 24 MASCO__Y6 $T=534265 146895 0 0 $X=534265 $Y=146895
X603 24 MASCO__Y6 $T=545265 50835 0 0 $X=545265 $Y=50835
X604 24 MASCO__Y6 $T=545265 146895 0 0 $X=545265 $Y=146895
X605 23 MASCO__Y7 $T=378695 51895 0 0 $X=378695 $Y=51895
X606 23 MASCO__Y7 $T=378695 56895 0 0 $X=378695 $Y=56895
X607 23 MASCO__Y7 $T=378695 61895 0 0 $X=378695 $Y=61895
X608 23 MASCO__Y7 $T=378695 66895 0 0 $X=378695 $Y=66895
X609 23 MASCO__Y7 $T=378695 71895 0 0 $X=378695 $Y=71895
X610 23 MASCO__Y7 $T=378695 76895 0 0 $X=378695 $Y=76895
X611 23 MASCO__Y7 $T=378695 81895 0 0 $X=378695 $Y=81895
X612 23 MASCO__Y7 $T=378695 86895 0 0 $X=378695 $Y=86895
X613 23 MASCO__Y7 $T=378695 91895 0 0 $X=378695 $Y=91895
X614 23 MASCO__Y7 $T=378695 96895 0 0 $X=378695 $Y=96895
X615 23 MASCO__Y7 $T=378695 101895 0 0 $X=378695 $Y=101895
X616 23 MASCO__Y7 $T=378695 106895 0 0 $X=378695 $Y=106895
X617 23 MASCO__Y7 $T=378695 111895 0 0 $X=378695 $Y=111895
X618 23 MASCO__Y7 $T=378695 116895 0 0 $X=378695 $Y=116895
X619 23 MASCO__Y7 $T=378695 121895 0 0 $X=378695 $Y=121895
X620 23 MASCO__Y7 $T=378695 126895 0 0 $X=378695 $Y=126895
X621 23 MASCO__Y7 $T=378695 131895 0 0 $X=378695 $Y=131895
X622 23 MASCO__Y7 $T=378695 136895 0 0 $X=378695 $Y=136895
X623 23 MASCO__Y7 $T=378695 141895 0 0 $X=378695 $Y=141895
X624 23 MASCO__Y7 $T=396695 51895 0 0 $X=396695 $Y=51895
X625 23 MASCO__Y7 $T=396695 56895 0 0 $X=396695 $Y=56895
X626 23 MASCO__Y7 $T=396695 61895 0 0 $X=396695 $Y=61895
X627 23 MASCO__Y7 $T=396695 66895 0 0 $X=396695 $Y=66895
X628 23 MASCO__Y7 $T=396695 71895 0 0 $X=396695 $Y=71895
X629 23 MASCO__Y7 $T=396695 76895 0 0 $X=396695 $Y=76895
X630 23 MASCO__Y7 $T=396695 81895 0 0 $X=396695 $Y=81895
X631 23 MASCO__Y7 $T=396695 86895 0 0 $X=396695 $Y=86895
X632 23 MASCO__Y7 $T=396695 91895 0 0 $X=396695 $Y=91895
X633 23 MASCO__Y7 $T=396695 96895 0 0 $X=396695 $Y=96895
X634 23 MASCO__Y7 $T=396695 101895 0 0 $X=396695 $Y=101895
X635 23 MASCO__Y7 $T=396695 106895 0 0 $X=396695 $Y=106895
X636 23 MASCO__Y7 $T=396695 111895 0 0 $X=396695 $Y=111895
X637 23 MASCO__Y7 $T=396695 116895 0 0 $X=396695 $Y=116895
X638 23 MASCO__Y7 $T=396695 121895 0 0 $X=396695 $Y=121895
X639 23 MASCO__Y7 $T=396695 126895 0 0 $X=396695 $Y=126895
X640 23 MASCO__Y7 $T=396695 131895 0 0 $X=396695 $Y=131895
X641 23 MASCO__Y7 $T=396695 136895 0 0 $X=396695 $Y=136895
X642 23 MASCO__Y7 $T=396695 141895 0 0 $X=396695 $Y=141895
X643 23 MASCO__Y7 $T=414695 51895 0 0 $X=414695 $Y=51895
X644 23 MASCO__Y7 $T=414695 56895 0 0 $X=414695 $Y=56895
X645 23 MASCO__Y7 $T=414695 61895 0 0 $X=414695 $Y=61895
X646 23 MASCO__Y7 $T=414695 66895 0 0 $X=414695 $Y=66895
X647 23 MASCO__Y7 $T=414695 71895 0 0 $X=414695 $Y=71895
X648 23 MASCO__Y7 $T=414695 76895 0 0 $X=414695 $Y=76895
X649 23 MASCO__Y7 $T=414695 81895 0 0 $X=414695 $Y=81895
X650 23 MASCO__Y7 $T=414695 86895 0 0 $X=414695 $Y=86895
X651 23 MASCO__Y7 $T=414695 91895 0 0 $X=414695 $Y=91895
X652 23 MASCO__Y7 $T=414695 96895 0 0 $X=414695 $Y=96895
X653 23 MASCO__Y7 $T=414695 101895 0 0 $X=414695 $Y=101895
X654 23 MASCO__Y7 $T=414695 106895 0 0 $X=414695 $Y=106895
X655 23 MASCO__Y7 $T=414695 111895 0 0 $X=414695 $Y=111895
X656 23 MASCO__Y7 $T=414695 116895 0 0 $X=414695 $Y=116895
X657 23 MASCO__Y7 $T=414695 121895 0 0 $X=414695 $Y=121895
X658 23 MASCO__Y7 $T=414695 126895 0 0 $X=414695 $Y=126895
X659 23 MASCO__Y7 $T=414695 131895 0 0 $X=414695 $Y=131895
X660 23 MASCO__Y7 $T=414695 136895 0 0 $X=414695 $Y=136895
X661 23 MASCO__Y7 $T=414695 141895 0 0 $X=414695 $Y=141895
X662 24 MASCO__Y7 $T=502265 51895 0 0 $X=502265 $Y=51895
X663 24 MASCO__Y7 $T=502265 56895 0 0 $X=502265 $Y=56895
X664 24 MASCO__Y7 $T=502265 61895 0 0 $X=502265 $Y=61895
X665 24 MASCO__Y7 $T=502265 66895 0 0 $X=502265 $Y=66895
X666 24 MASCO__Y7 $T=502265 71895 0 0 $X=502265 $Y=71895
X667 24 MASCO__Y7 $T=502265 76895 0 0 $X=502265 $Y=76895
X668 24 MASCO__Y7 $T=502265 81895 0 0 $X=502265 $Y=81895
X669 24 MASCO__Y7 $T=502265 86895 0 0 $X=502265 $Y=86895
X670 24 MASCO__Y7 $T=502265 91895 0 0 $X=502265 $Y=91895
X671 24 MASCO__Y7 $T=502265 96895 0 0 $X=502265 $Y=96895
X672 24 MASCO__Y7 $T=502265 101895 0 0 $X=502265 $Y=101895
X673 24 MASCO__Y7 $T=502265 106895 0 0 $X=502265 $Y=106895
X674 24 MASCO__Y7 $T=502265 111895 0 0 $X=502265 $Y=111895
X675 24 MASCO__Y7 $T=502265 116895 0 0 $X=502265 $Y=116895
X676 24 MASCO__Y7 $T=502265 121895 0 0 $X=502265 $Y=121895
X677 24 MASCO__Y7 $T=502265 126895 0 0 $X=502265 $Y=126895
X678 24 MASCO__Y7 $T=502265 131895 0 0 $X=502265 $Y=131895
X679 24 MASCO__Y7 $T=502265 136895 0 0 $X=502265 $Y=136895
X680 24 MASCO__Y7 $T=502265 141895 0 0 $X=502265 $Y=141895
X681 24 MASCO__Y7 $T=520265 51895 0 0 $X=520265 $Y=51895
X682 24 MASCO__Y7 $T=520265 56895 0 0 $X=520265 $Y=56895
X683 24 MASCO__Y7 $T=520265 61895 0 0 $X=520265 $Y=61895
X684 24 MASCO__Y7 $T=520265 66895 0 0 $X=520265 $Y=66895
X685 24 MASCO__Y7 $T=520265 71895 0 0 $X=520265 $Y=71895
X686 24 MASCO__Y7 $T=520265 76895 0 0 $X=520265 $Y=76895
X687 24 MASCO__Y7 $T=520265 81895 0 0 $X=520265 $Y=81895
X688 24 MASCO__Y7 $T=520265 86895 0 0 $X=520265 $Y=86895
X689 24 MASCO__Y7 $T=520265 91895 0 0 $X=520265 $Y=91895
X690 24 MASCO__Y7 $T=520265 96895 0 0 $X=520265 $Y=96895
X691 24 MASCO__Y7 $T=520265 101895 0 0 $X=520265 $Y=101895
X692 24 MASCO__Y7 $T=520265 106895 0 0 $X=520265 $Y=106895
X693 24 MASCO__Y7 $T=520265 111895 0 0 $X=520265 $Y=111895
X694 24 MASCO__Y7 $T=520265 116895 0 0 $X=520265 $Y=116895
X695 24 MASCO__Y7 $T=520265 121895 0 0 $X=520265 $Y=121895
X696 24 MASCO__Y7 $T=520265 126895 0 0 $X=520265 $Y=126895
X697 24 MASCO__Y7 $T=520265 131895 0 0 $X=520265 $Y=131895
X698 24 MASCO__Y7 $T=520265 136895 0 0 $X=520265 $Y=136895
X699 24 MASCO__Y7 $T=520265 141895 0 0 $X=520265 $Y=141895
X700 24 MASCO__Y7 $T=538265 51895 0 0 $X=538265 $Y=51895
X701 24 MASCO__Y7 $T=538265 56895 0 0 $X=538265 $Y=56895
X702 24 MASCO__Y7 $T=538265 61895 0 0 $X=538265 $Y=61895
X703 24 MASCO__Y7 $T=538265 66895 0 0 $X=538265 $Y=66895
X704 24 MASCO__Y7 $T=538265 71895 0 0 $X=538265 $Y=71895
X705 24 MASCO__Y7 $T=538265 76895 0 0 $X=538265 $Y=76895
X706 24 MASCO__Y7 $T=538265 81895 0 0 $X=538265 $Y=81895
X707 24 MASCO__Y7 $T=538265 86895 0 0 $X=538265 $Y=86895
X708 24 MASCO__Y7 $T=538265 91895 0 0 $X=538265 $Y=91895
X709 24 MASCO__Y7 $T=538265 96895 0 0 $X=538265 $Y=96895
X710 24 MASCO__Y7 $T=538265 101895 0 0 $X=538265 $Y=101895
X711 24 MASCO__Y7 $T=538265 106895 0 0 $X=538265 $Y=106895
X712 24 MASCO__Y7 $T=538265 111895 0 0 $X=538265 $Y=111895
X713 24 MASCO__Y7 $T=538265 116895 0 0 $X=538265 $Y=116895
X714 24 MASCO__Y7 $T=538265 121895 0 0 $X=538265 $Y=121895
X715 24 MASCO__Y7 $T=538265 126895 0 0 $X=538265 $Y=126895
X716 24 MASCO__Y7 $T=538265 131895 0 0 $X=538265 $Y=131895
X717 24 MASCO__Y7 $T=538265 136895 0 0 $X=538265 $Y=136895
X718 24 MASCO__Y7 $T=538265 141895 0 0 $X=538265 $Y=141895
X719 23 MASCO__Y8 $T=377695 52895 0 0 $X=377695 $Y=52895
X720 23 MASCO__Y8 $T=377695 76895 0 0 $X=377695 $Y=76895
X721 23 MASCO__Y8 $T=377695 100895 0 0 $X=377695 $Y=100895
X722 23 MASCO__Y8 $T=391695 52895 0 0 $X=391695 $Y=52895
X723 23 MASCO__Y8 $T=391695 76895 0 0 $X=391695 $Y=76895
X724 23 MASCO__Y8 $T=391695 100895 0 0 $X=391695 $Y=100895
X725 23 MASCO__Y8 $T=405695 52895 0 0 $X=405695 $Y=52895
X726 23 MASCO__Y8 $T=405695 76895 0 0 $X=405695 $Y=76895
X727 23 MASCO__Y8 $T=405695 100895 0 0 $X=405695 $Y=100895
X728 23 MASCO__Y8 $T=419695 52895 0 0 $X=419695 $Y=52895
X729 23 MASCO__Y8 $T=419695 76895 0 0 $X=419695 $Y=76895
X730 23 MASCO__Y8 $T=419695 100895 0 0 $X=419695 $Y=100895
X731 24 MASCO__Y8 $T=501265 52895 0 0 $X=501265 $Y=52895
X732 24 MASCO__Y8 $T=501265 76895 0 0 $X=501265 $Y=76895
X733 24 MASCO__Y8 $T=501265 100895 0 0 $X=501265 $Y=100895
X734 24 MASCO__Y8 $T=515265 52895 0 0 $X=515265 $Y=52895
X735 24 MASCO__Y8 $T=515265 76895 0 0 $X=515265 $Y=76895
X736 24 MASCO__Y8 $T=515265 100895 0 0 $X=515265 $Y=100895
X737 24 MASCO__Y8 $T=529265 52895 0 0 $X=529265 $Y=52895
X738 24 MASCO__Y8 $T=529265 76895 0 0 $X=529265 $Y=76895
X739 24 MASCO__Y8 $T=529265 100895 0 0 $X=529265 $Y=100895
X740 24 MASCO__Y8 $T=543265 52895 0 0 $X=543265 $Y=52895
X741 24 MASCO__Y8 $T=543265 76895 0 0 $X=543265 $Y=76895
X742 24 MASCO__Y8 $T=543265 100895 0 0 $X=543265 $Y=100895
X743 23 MASCO__Y9 $T=377695 124895 0 0 $X=377695 $Y=124895
X744 23 MASCO__Y9 $T=391695 124895 0 0 $X=391695 $Y=124895
X745 23 MASCO__Y9 $T=405695 124895 0 0 $X=405695 $Y=124895
X746 23 MASCO__Y9 $T=419695 124895 0 0 $X=419695 $Y=124895
X747 24 MASCO__Y9 $T=501265 124895 0 0 $X=501265 $Y=124895
X748 24 MASCO__Y9 $T=515265 124895 0 0 $X=515265 $Y=124895
X749 24 MASCO__Y9 $T=529265 124895 0 0 $X=529265 $Y=124895
X750 24 MASCO__Y9 $T=543265 124895 0 0 $X=543265 $Y=124895
X751 14 9 9 MOSVC3 w=2e-05 l=3e-05 $X=16180 $Y=110530 $dt=3
X752 14 9 9 MOSVC3 w=2e-05 l=3e-05 $X=16180 $Y=132530 $dt=3
X753 14 9 9 MOSVC3 w=2e-05 l=3e-05 $X=48780 $Y=110530 $dt=3
X754 14 9 9 MOSVC3 w=2e-05 l=3e-05 $X=48780 $Y=132530 $dt=3
R4 9 25 5 $[s_res] $X=263280 $Y=3815 $dt=4
D5 9 14 p_dnw AREA=3.57048e-11 PJ=3.588e-05 perimeter=3.588e-05 $X=11740 $Y=84695 $dt=5
D6 9 14 p_dnw AREA=1.90124e-10 PJ=7.516e-05 perimeter=7.516e-05 $X=59815 $Y=81480 $dt=5
D7 9 14 p_dnw AREA=1.58288e-09 PJ=0.00049318 perimeter=0.00049318 $X=99710 $Y=59910 $dt=5
D8 9 14 p_dnw AREA=3.09086e-09 PJ=0.00032604 perimeter=0.00032604 $X=101390 $Y=114415 $dt=5
D9 9 7 p_dnw AREA=1.82058e-10 PJ=5.826e-05 perimeter=5.826e-05 $X=105905 $Y=15300 $dt=5
D10 9 8 p_dnw AREA=1.82058e-10 PJ=5.826e-05 perimeter=5.826e-05 $X=105905 $Y=44920 $dt=5
D11 9 8 p_dnw AREA=1.82058e-10 PJ=5.826e-05 perimeter=5.826e-05 $X=160185 $Y=15300 $dt=5
D12 9 7 p_dnw AREA=1.82058e-10 PJ=5.826e-05 perimeter=5.826e-05 $X=160185 $Y=44920 $dt=5
D13 9 14 p_dnw AREA=8.36476e-09 PJ=0.0003905 perimeter=0.0003905 $X=226790 $Y=95600 $dt=5
D14 9 14 p_dnw3 AREA=4.20992e-11 PJ=0 perimeter=0 $X=12880 $Y=85835 $dt=6
D15 9 9 p_dnw3 AREA=5.9176e-11 PJ=0.00010492 perimeter=0.00010492 $X=15380 $Y=110100 $dt=6
D16 9 9 p_dnw3 AREA=5.9176e-11 PJ=0.00010492 perimeter=0.00010492 $X=15380 $Y=132100 $dt=6
D17 9 9 p_dnw3 AREA=5.9176e-11 PJ=0.00010492 perimeter=0.00010492 $X=47980 $Y=110100 $dt=6
D18 9 9 p_dnw3 AREA=5.9176e-11 PJ=0.00010492 perimeter=0.00010492 $X=47980 $Y=132100 $dt=6
D19 9 14 p_dnw3 AREA=1.56539e-10 PJ=0 perimeter=0 $X=61455 $Y=83900 $dt=6
D20 9 7 p_dnw3 AREA=5.86064e-10 PJ=7.406e-05 perimeter=7.406e-05 $X=105905 $Y=18860 $dt=6
D21 9 8 p_dnw3 AREA=5.86064e-10 PJ=7.406e-05 perimeter=7.406e-05 $X=105905 $Y=33460 $dt=6
D22 9 14 p_dnw3 AREA=1.22554e-09 PJ=0 perimeter=0 $X=108190 $Y=68670 $dt=6
D23 9 14 p_dnw3 AREA=1.15225e-09 PJ=0.00012214 perimeter=0.00012214 $X=108190 $Y=82290 $dt=6
D24 9 14 p_dnw3 AREA=1.15028e-09 PJ=0 perimeter=0 $X=112150 $Y=124955 $dt=6
D25 9 14 p_dnw3 AREA=1.15028e-09 PJ=0 perimeter=0 $X=112150 $Y=137935 $dt=6
D26 9 8 p_dnw3 AREA=5.86064e-10 PJ=7.406e-05 perimeter=7.406e-05 $X=160185 $Y=18860 $dt=6
D27 9 7 p_dnw3 AREA=5.86064e-10 PJ=7.406e-05 perimeter=7.406e-05 $X=160185 $Y=33460 $dt=6
C28 11 26 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=231620 $Y=128940 $dt=9
C29 11 26 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=263220 $Y=97740 $dt=9
C30 11 26 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=263220 $Y=128940 $dt=9
C31 11 26 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=294820 $Y=97740 $dt=9
C32 11 26 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=294820 $Y=128940 $dt=9
C33 11 26 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=326420 $Y=97740 $dt=9
C34 11 26 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=326420 $Y=128940 $dt=9
.ends current_source_gm_10_en_r
