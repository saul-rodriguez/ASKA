* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : bandgap_su                                   *
* Netlisted  : Mon Aug 26 08:15:29 2024                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(ne3) nem ndiff(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 1 MP(pe3) pem pdiff(D) p1trm(G) pdiff(S) nwtrm(B)
*.DEVTMPLT 2 Q(qpvc3) qpvmc bulk(C) nwtrm(B) pdiff(E)
*.DEVTMPLT 3 D(p_dnw) p_dnw bulk(POS) nwtrm(NEG)
*.DEVTMPLT 4 D(p_dnw3) p_dnwm bulk(POS) nwtrm(NEG)
*.DEVTMPLT 5 R(rpp1k1_3) rpp1k1_s p1trm(POS) p1trm(NEG) bulk(SUB)
*.DEVTMPLT 6 C(cmm5t) cmim capm(POS) m4trm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724652923740                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724652923740 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724652923740

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_724652923741                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_724652923741 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_724652923741

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724652923742                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724652923742 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724652923742

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_724652923743                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_724652923743 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_724652923743

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_724652923744                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_724652923744 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_724652923744

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724652923745                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724652923745 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724652923745

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724652923746                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724652923746 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724652923746

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724652923748                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724652923748 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724652923748

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_724652923749                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_724652923749 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_724652923749

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246529237410                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246529237410 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246529237410

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246529237412                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246529237412 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246529237412

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246529237414                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246529237414 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246529237414

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246529237415                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246529237415 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246529237415

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246529237420                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246529237420 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246529237420

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246529237422                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246529237422 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246529237422

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246529237424                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246529237424 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246529237424

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246529237429                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246529237429 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246529237429

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724652923740                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724652923740 1 2 3 4 5
** N=5 EP=5 FDC=5
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=1
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=1
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=1
D4 5 4 p_dnw3 AREA=1.04198e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=4
.ends pe3_CDNS_724652923740

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724652923741                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724652923741 1 2 3 4
** N=4 EP=4 FDC=4
M0 3 2 1 4 ne3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
M1 1 2 3 4 ne3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=0
M2 3 2 1 4 ne3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=0
M3 1 2 3 4 ne3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=0
.ends ne3_CDNS_724652923741

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_724652923742                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_724652923742 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.0005215 W=8e-06 $[rpp1k1_3] $SUB=3 $X=-8220 $Y=0 $dt=5
.ends rpp1k1_3_CDNS_724652923742

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_724652923743                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_724652923743 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.00082283 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=5
.ends rpp1k1_3_CDNS_724652923743

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724652923744                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724652923744 1 2 3 4
** N=4 EP=4 FDC=1
M0 3 2 1 4 ne3 L=1e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
.ends ne3_CDNS_724652923744

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724652923746                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724652923746 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=1
M0 3 2 1 4 pe3 L=5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_724652923746

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724652923747                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724652923747 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 3 2 1 4 pe3 L=5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
D1 5 4 p_dnw3 AREA=9.67212e-11 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=4
.ends pe3_CDNS_724652923747

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724652923748                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724652923748 1 2 3
** N=3 EP=3 FDC=1
M0 2 2 1 3 ne3 L=2e-06 W=1e-06 AD=4.8e-13 AS=4.8e-13 PD=2.96e-06 PS=2.96e-06 $X=0 $Y=0 $dt=0
.ends ne3_CDNS_724652923748

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724652923749                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724652923749 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
M0 3 2 1 1 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_724652923749

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7246529237410                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7246529237410 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
.ends ne3_CDNS_7246529237410

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7246529237411                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7246529237411 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.00082283 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=5
.ends rpp1k1_3_CDNS_7246529237411

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: bandgap_su                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt bandgap_su 5 6 7 3
** N=24 EP=4 FDC=165
X0 1 VIA1_C_CDNS_724652923740 $T=9365 74485 0 0 $X=9225 $Y=73775
X1 2 VIA1_C_CDNS_724652923740 $T=10075 52335 0 0 $X=9935 $Y=51625
X2 3 VIA1_C_CDNS_724652923740 $T=10390 104220 0 0 $X=10250 $Y=103510
X3 3 VIA1_C_CDNS_724652923740 $T=10390 131040 0 0 $X=10250 $Y=130330
X4 4 VIA1_C_CDNS_724652923740 $T=10905 76265 0 0 $X=10765 $Y=75555
X5 5 VIA1_C_CDNS_724652923740 $T=11615 54115 0 0 $X=11475 $Y=53405
X6 3 VIA1_C_CDNS_724652923740 $T=11930 104220 0 0 $X=11790 $Y=103510
X7 3 VIA1_C_CDNS_724652923740 $T=11930 131040 0 0 $X=11790 $Y=130330
X8 1 VIA1_C_CDNS_724652923740 $T=12445 74485 0 0 $X=12305 $Y=73775
X9 3 VIA1_C_CDNS_724652923740 $T=12630 104220 0 0 $X=12490 $Y=103510
X10 3 VIA1_C_CDNS_724652923740 $T=12630 131040 0 0 $X=12490 $Y=130330
X11 6 VIA1_C_CDNS_724652923740 $T=12860 15465 0 0 $X=12720 $Y=14755
X12 6 VIA1_C_CDNS_724652923740 $T=12860 40105 0 0 $X=12720 $Y=39395
X13 2 VIA1_C_CDNS_724652923740 $T=13155 52335 0 0 $X=13015 $Y=51625
X14 4 VIA1_C_CDNS_724652923740 $T=13985 76265 0 0 $X=13845 $Y=75555
X15 7 VIA1_C_CDNS_724652923740 $T=14170 98880 0 0 $X=14030 $Y=98170
X16 7 VIA1_C_CDNS_724652923740 $T=14170 132820 0 0 $X=14030 $Y=132110
X17 6 VIA1_C_CDNS_724652923740 $T=14400 15465 0 0 $X=14260 $Y=14755
X18 6 VIA1_C_CDNS_724652923740 $T=14400 40105 0 0 $X=14260 $Y=39395
X19 5 VIA1_C_CDNS_724652923740 $T=14695 54115 0 0 $X=14555 $Y=53405
X20 3 VIA1_C_CDNS_724652923740 $T=14870 104220 0 0 $X=14730 $Y=103510
X21 3 VIA1_C_CDNS_724652923740 $T=14870 131040 0 0 $X=14730 $Y=130330
X22 6 VIA1_C_CDNS_724652923740 $T=15100 15465 0 0 $X=14960 $Y=14755
X23 6 VIA1_C_CDNS_724652923740 $T=15100 40105 0 0 $X=14960 $Y=39395
X24 1 VIA1_C_CDNS_724652923740 $T=15525 74485 0 0 $X=15385 $Y=73775
X25 2 VIA1_C_CDNS_724652923740 $T=16235 52335 0 0 $X=16095 $Y=51625
X26 7 VIA1_C_CDNS_724652923740 $T=16410 98880 0 0 $X=16270 $Y=98170
X27 7 VIA1_C_CDNS_724652923740 $T=16410 132820 0 0 $X=16270 $Y=132110
X28 8 VIA1_C_CDNS_724652923740 $T=16640 11905 0 0 $X=16500 $Y=11195
X29 2 VIA1_C_CDNS_724652923740 $T=16640 43665 0 0 $X=16500 $Y=42955
X30 3 VIA1_C_CDNS_724652923740 $T=17110 104220 0 0 $X=16970 $Y=103510
X31 3 VIA1_C_CDNS_724652923740 $T=17110 131040 0 0 $X=16970 $Y=130330
X32 6 VIA1_C_CDNS_724652923740 $T=17340 15465 0 0 $X=17200 $Y=14755
X33 6 VIA1_C_CDNS_724652923740 $T=17340 40105 0 0 $X=17200 $Y=39395
X34 9 VIA1_C_CDNS_724652923740 $T=18650 102440 0 0 $X=18510 $Y=101730
X35 1 VIA1_C_CDNS_724652923740 $T=18650 134600 0 0 $X=18510 $Y=133890
X36 2 VIA1_C_CDNS_724652923740 $T=18880 13685 0 0 $X=18740 $Y=12975
X37 8 VIA1_C_CDNS_724652923740 $T=18880 41885 0 0 $X=18740 $Y=41175
X38 3 VIA1_C_CDNS_724652923740 $T=19350 104220 0 0 $X=19210 $Y=103510
X39 3 VIA1_C_CDNS_724652923740 $T=19350 131040 0 0 $X=19210 $Y=130330
X40 6 VIA1_C_CDNS_724652923740 $T=19580 15465 0 0 $X=19440 $Y=14755
X41 6 VIA1_C_CDNS_724652923740 $T=19580 40105 0 0 $X=19440 $Y=39395
X42 7 VIA1_C_CDNS_724652923740 $T=20890 98880 0 0 $X=20750 $Y=98170
X43 7 VIA1_C_CDNS_724652923740 $T=20890 132820 0 0 $X=20750 $Y=132110
X44 10 VIA1_C_CDNS_724652923740 $T=21120 10125 0 0 $X=20980 $Y=9415
X45 11 VIA1_C_CDNS_724652923740 $T=21120 45445 0 0 $X=20980 $Y=44735
X46 3 VIA1_C_CDNS_724652923740 $T=21590 104220 0 0 $X=21450 $Y=103510
X47 3 VIA1_C_CDNS_724652923740 $T=21590 131040 0 0 $X=21450 $Y=130330
X48 6 VIA1_C_CDNS_724652923740 $T=21820 15465 0 0 $X=21680 $Y=14755
X49 6 VIA1_C_CDNS_724652923740 $T=21820 40105 0 0 $X=21680 $Y=39395
X50 8 VIA1_C_CDNS_724652923740 $T=22460 54255 0 0 $X=22320 $Y=53545
X51 7 VIA1_C_CDNS_724652923740 $T=23130 98880 0 0 $X=22990 $Y=98170
X52 7 VIA1_C_CDNS_724652923740 $T=23130 132820 0 0 $X=22990 $Y=132110
X53 9 VIA1_C_CDNS_724652923740 $T=23170 76265 0 0 $X=23030 $Y=75555
X54 8 VIA1_C_CDNS_724652923740 $T=23360 11905 0 0 $X=23220 $Y=11195
X55 2 VIA1_C_CDNS_724652923740 $T=23360 43665 0 0 $X=23220 $Y=42955
X56 3 VIA1_C_CDNS_724652923740 $T=23830 104220 0 0 $X=23690 $Y=103510
X57 3 VIA1_C_CDNS_724652923740 $T=23830 131040 0 0 $X=23690 $Y=130330
X58 4 VIA1_C_CDNS_724652923740 $T=24000 52475 0 0 $X=23860 $Y=51765
X59 6 VIA1_C_CDNS_724652923740 $T=24060 15465 0 0 $X=23920 $Y=14755
X60 6 VIA1_C_CDNS_724652923740 $T=24060 40105 0 0 $X=23920 $Y=39395
X61 12 VIA1_C_CDNS_724652923740 $T=24710 74485 0 0 $X=24570 $Y=73775
X62 1 VIA1_C_CDNS_724652923740 $T=25370 100660 0 0 $X=25230 $Y=99950
X63 9 VIA1_C_CDNS_724652923740 $T=25370 136380 0 0 $X=25230 $Y=135670
X64 8 VIA1_C_CDNS_724652923740 $T=25540 54255 0 0 $X=25400 $Y=53545
X65 2 VIA1_C_CDNS_724652923740 $T=25600 13685 0 0 $X=25460 $Y=12975
X66 8 VIA1_C_CDNS_724652923740 $T=25600 41885 0 0 $X=25460 $Y=41175
X67 3 VIA1_C_CDNS_724652923740 $T=26070 104220 0 0 $X=25930 $Y=103510
X68 3 VIA1_C_CDNS_724652923740 $T=26070 131040 0 0 $X=25930 $Y=130330
X69 9 VIA1_C_CDNS_724652923740 $T=26250 76265 0 0 $X=26110 $Y=75555
X70 6 VIA1_C_CDNS_724652923740 $T=26300 15465 0 0 $X=26160 $Y=14755
X71 6 VIA1_C_CDNS_724652923740 $T=26300 40105 0 0 $X=26160 $Y=39395
X72 4 VIA1_C_CDNS_724652923740 $T=27080 52475 0 0 $X=26940 $Y=51765
X73 9 VIA1_C_CDNS_724652923740 $T=27610 102440 0 0 $X=27470 $Y=101730
X74 1 VIA1_C_CDNS_724652923740 $T=27610 134600 0 0 $X=27470 $Y=133890
X75 12 VIA1_C_CDNS_724652923740 $T=27790 74485 0 0 $X=27650 $Y=73775
X76 6 VIA1_C_CDNS_724652923740 $T=27840 15465 0 0 $X=27700 $Y=14755
X77 6 VIA1_C_CDNS_724652923740 $T=27840 40105 0 0 $X=27700 $Y=39395
X78 3 VIA1_C_CDNS_724652923740 $T=28310 104220 0 0 $X=28170 $Y=103510
X79 3 VIA1_C_CDNS_724652923740 $T=28310 131040 0 0 $X=28170 $Y=130330
X80 8 VIA1_C_CDNS_724652923740 $T=28620 54255 0 0 $X=28480 $Y=53545
X81 9 VIA1_C_CDNS_724652923740 $T=29330 76265 0 0 $X=29190 $Y=75555
X82 7 VIA1_C_CDNS_724652923740 $T=29850 98880 0 0 $X=29710 $Y=98170
X83 7 VIA1_C_CDNS_724652923740 $T=29850 132820 0 0 $X=29710 $Y=132110
X84 3 VIA1_C_CDNS_724652923740 $T=30550 104220 0 0 $X=30410 $Y=103510
X85 3 VIA1_C_CDNS_724652923740 $T=30550 131040 0 0 $X=30410 $Y=130330
X86 7 VIA1_C_CDNS_724652923740 $T=32090 98880 0 0 $X=31950 $Y=98170
X87 7 VIA1_C_CDNS_724652923740 $T=32090 132820 0 0 $X=31950 $Y=132110
X88 3 VIA1_C_CDNS_724652923740 $T=32790 104220 0 0 $X=32650 $Y=103510
X89 3 VIA1_C_CDNS_724652923740 $T=32790 131040 0 0 $X=32650 $Y=130330
X90 1 VIA1_C_CDNS_724652923740 $T=34330 100660 0 0 $X=34190 $Y=99950
X91 9 VIA1_C_CDNS_724652923740 $T=34330 136380 0 0 $X=34190 $Y=135670
X92 3 VIA1_C_CDNS_724652923740 $T=35030 104220 0 0 $X=34890 $Y=103510
X93 3 VIA1_C_CDNS_724652923740 $T=35030 131040 0 0 $X=34890 $Y=130330
X94 7 VIA1_C_CDNS_724652923740 $T=36570 98880 0 0 $X=36430 $Y=98170
X95 7 VIA1_C_CDNS_724652923740 $T=36570 132820 0 0 $X=36430 $Y=132110
X96 3 VIA1_C_CDNS_724652923740 $T=37270 104220 0 0 $X=37130 $Y=103510
X97 3 VIA1_C_CDNS_724652923740 $T=37270 131040 0 0 $X=37130 $Y=130330
X98 7 VIA1_C_CDNS_724652923740 $T=38810 98880 0 0 $X=38670 $Y=98170
X99 7 VIA1_C_CDNS_724652923740 $T=38810 132820 0 0 $X=38670 $Y=132110
X100 3 VIA1_C_CDNS_724652923740 $T=39510 104220 0 0 $X=39370 $Y=103510
X101 3 VIA1_C_CDNS_724652923740 $T=39510 131040 0 0 $X=39370 $Y=130330
X102 3 VIA1_C_CDNS_724652923740 $T=41050 104220 0 0 $X=40910 $Y=103510
X103 3 VIA1_C_CDNS_724652923740 $T=41050 131040 0 0 $X=40910 $Y=130330
X104 12 VIA1_C_CDNS_724652923740 $T=42835 58225 0 0 $X=42695 $Y=57515
X105 12 VIA1_C_CDNS_724652923740 $T=42835 85685 0 0 $X=42695 $Y=84975
X106 6 VIA1_C_CDNS_724652923740 $T=44510 14010 0 0 $X=44370 $Y=13300
X107 6 VIA1_C_CDNS_724652923740 $T=44510 38730 0 0 $X=44370 $Y=38020
X108 12 VIA1_C_CDNS_724652923740 $T=48375 58225 0 0 $X=48235 $Y=57515
X109 12 VIA1_C_CDNS_724652923740 $T=48375 85685 0 0 $X=48235 $Y=84975
X110 12 VIA1_C_CDNS_724652923740 $T=49075 58225 0 0 $X=48935 $Y=57515
X111 12 VIA1_C_CDNS_724652923740 $T=49075 85685 0 0 $X=48935 $Y=84975
X112 6 VIA1_C_CDNS_724652923740 $T=50050 14010 0 0 $X=49910 $Y=13300
X113 6 VIA1_C_CDNS_724652923740 $T=50050 38730 0 0 $X=49910 $Y=38020
X114 6 VIA1_C_CDNS_724652923740 $T=50750 14010 0 0 $X=50610 $Y=13300
X115 6 VIA1_C_CDNS_724652923740 $T=50750 38730 0 0 $X=50610 $Y=38020
X116 13 VIA1_C_CDNS_724652923740 $T=54615 54665 0 0 $X=54475 $Y=53955
X117 14 VIA1_C_CDNS_724652923740 $T=54615 89245 0 0 $X=54475 $Y=88535
X118 12 VIA1_C_CDNS_724652923740 $T=55315 58225 0 0 $X=55175 $Y=57515
X119 12 VIA1_C_CDNS_724652923740 $T=55315 85685 0 0 $X=55175 $Y=84975
X120 14 VIA1_C_CDNS_724652923740 $T=56290 12230 0 0 $X=56150 $Y=11520
X121 13 VIA1_C_CDNS_724652923740 $T=56290 40510 0 0 $X=56150 $Y=39800
X122 6 VIA1_C_CDNS_724652923740 $T=56990 14010 0 0 $X=56850 $Y=13300
X123 6 VIA1_C_CDNS_724652923740 $T=56990 38730 0 0 $X=56850 $Y=38020
X124 14 VIA1_C_CDNS_724652923740 $T=60855 56445 0 0 $X=60715 $Y=55735
X125 13 VIA1_C_CDNS_724652923740 $T=60855 87465 0 0 $X=60715 $Y=86755
X126 12 VIA1_C_CDNS_724652923740 $T=61555 58225 0 0 $X=61415 $Y=57515
X127 12 VIA1_C_CDNS_724652923740 $T=61555 85685 0 0 $X=61415 $Y=84975
X128 13 VIA1_C_CDNS_724652923740 $T=62530 10450 0 0 $X=62390 $Y=9740
X129 14 VIA1_C_CDNS_724652923740 $T=62530 42290 0 0 $X=62390 $Y=41580
X130 6 VIA1_C_CDNS_724652923740 $T=63230 14010 0 0 $X=63090 $Y=13300
X131 6 VIA1_C_CDNS_724652923740 $T=63230 38730 0 0 $X=63090 $Y=38020
X132 13 VIA1_C_CDNS_724652923740 $T=67095 54665 0 0 $X=66955 $Y=53955
X133 14 VIA1_C_CDNS_724652923740 $T=67095 89245 0 0 $X=66955 $Y=88535
X134 12 VIA1_C_CDNS_724652923740 $T=67795 58225 0 0 $X=67655 $Y=57515
X135 12 VIA1_C_CDNS_724652923740 $T=67795 85685 0 0 $X=67655 $Y=84975
X136 14 VIA1_C_CDNS_724652923740 $T=68770 12230 0 0 $X=68630 $Y=11520
X137 13 VIA1_C_CDNS_724652923740 $T=68770 40510 0 0 $X=68630 $Y=39800
X138 6 VIA1_C_CDNS_724652923740 $T=69470 14010 0 0 $X=69330 $Y=13300
X139 6 VIA1_C_CDNS_724652923740 $T=69470 38730 0 0 $X=69330 $Y=38020
X140 14 VIA1_C_CDNS_724652923740 $T=73335 56445 0 0 $X=73195 $Y=55735
X141 13 VIA1_C_CDNS_724652923740 $T=73335 87465 0 0 $X=73195 $Y=86755
X142 12 VIA1_C_CDNS_724652923740 $T=74035 58225 0 0 $X=73895 $Y=57515
X143 12 VIA1_C_CDNS_724652923740 $T=74035 85685 0 0 $X=73895 $Y=84975
X144 13 VIA1_C_CDNS_724652923740 $T=75010 10450 0 0 $X=74870 $Y=9740
X145 14 VIA1_C_CDNS_724652923740 $T=75010 42290 0 0 $X=74870 $Y=41580
X146 6 VIA1_C_CDNS_724652923740 $T=75710 14010 0 0 $X=75570 $Y=13300
X147 6 VIA1_C_CDNS_724652923740 $T=75710 38730 0 0 $X=75570 $Y=38020
X148 3 VIA1_C_CDNS_724652923740 $T=78805 123400 0 0 $X=78665 $Y=122690
X149 13 VIA1_C_CDNS_724652923740 $T=79575 54665 0 0 $X=79435 $Y=53955
X150 14 VIA1_C_CDNS_724652923740 $T=79575 89245 0 0 $X=79435 $Y=88535
X151 12 VIA1_C_CDNS_724652923740 $T=80275 58225 0 0 $X=80135 $Y=57515
X152 12 VIA1_C_CDNS_724652923740 $T=80275 85685 0 0 $X=80135 $Y=84975
X153 14 VIA1_C_CDNS_724652923740 $T=81250 12230 0 0 $X=81110 $Y=11520
X154 13 VIA1_C_CDNS_724652923740 $T=81250 40510 0 0 $X=81110 $Y=39800
X155 6 VIA1_C_CDNS_724652923740 $T=81950 14010 0 0 $X=81810 $Y=13300
X156 6 VIA1_C_CDNS_724652923740 $T=81950 38730 0 0 $X=81810 $Y=38020
X157 15 VIA1_C_CDNS_724652923740 $T=84345 121620 0 0 $X=84205 $Y=120910
X158 3 VIA1_C_CDNS_724652923740 $T=85045 123400 0 0 $X=84905 $Y=122690
X159 14 VIA1_C_CDNS_724652923740 $T=85815 56445 0 0 $X=85675 $Y=55735
X160 13 VIA1_C_CDNS_724652923740 $T=85815 87465 0 0 $X=85675 $Y=86755
X161 12 VIA1_C_CDNS_724652923740 $T=86515 58225 0 0 $X=86375 $Y=57515
X162 12 VIA1_C_CDNS_724652923740 $T=86515 85685 0 0 $X=86375 $Y=84975
X163 13 VIA1_C_CDNS_724652923740 $T=87490 10450 0 0 $X=87350 $Y=9740
X164 14 VIA1_C_CDNS_724652923740 $T=87490 42290 0 0 $X=87350 $Y=41580
X165 6 VIA1_C_CDNS_724652923740 $T=88190 14010 0 0 $X=88050 $Y=13300
X166 6 VIA1_C_CDNS_724652923740 $T=88190 38730 0 0 $X=88050 $Y=38020
X167 16 VIA1_C_CDNS_724652923740 $T=90585 119840 0 0 $X=90445 $Y=119130
X168 13 VIA1_C_CDNS_724652923740 $T=92055 54665 0 0 $X=91915 $Y=53955
X169 14 VIA1_C_CDNS_724652923740 $T=92055 89245 0 0 $X=91915 $Y=88535
X170 12 VIA1_C_CDNS_724652923740 $T=92755 58225 0 0 $X=92615 $Y=57515
X171 12 VIA1_C_CDNS_724652923740 $T=92755 85685 0 0 $X=92615 $Y=84975
X172 14 VIA1_C_CDNS_724652923740 $T=93730 12230 0 0 $X=93590 $Y=11520
X173 13 VIA1_C_CDNS_724652923740 $T=93730 40510 0 0 $X=93590 $Y=39800
X174 6 VIA1_C_CDNS_724652923740 $T=94430 14010 0 0 $X=94290 $Y=13300
X175 6 VIA1_C_CDNS_724652923740 $T=94430 38730 0 0 $X=94290 $Y=38020
X176 14 VIA1_C_CDNS_724652923740 $T=98295 56445 0 0 $X=98155 $Y=55735
X177 13 VIA1_C_CDNS_724652923740 $T=98295 87465 0 0 $X=98155 $Y=86755
X178 12 VIA1_C_CDNS_724652923740 $T=98995 58225 0 0 $X=98855 $Y=57515
X179 12 VIA1_C_CDNS_724652923740 $T=98995 85685 0 0 $X=98855 $Y=84975
X180 13 VIA1_C_CDNS_724652923740 $T=99970 10450 0 0 $X=99830 $Y=9740
X181 14 VIA1_C_CDNS_724652923740 $T=99970 42290 0 0 $X=99830 $Y=41580
X182 6 VIA1_C_CDNS_724652923740 $T=100670 14010 0 0 $X=100530 $Y=13300
X183 6 VIA1_C_CDNS_724652923740 $T=100670 38730 0 0 $X=100530 $Y=38020
X184 12 VIA1_C_CDNS_724652923740 $T=104535 58225 0 0 $X=104395 $Y=57515
X185 12 VIA1_C_CDNS_724652923740 $T=104535 85685 0 0 $X=104395 $Y=84975
X186 6 VIA1_C_CDNS_724652923740 $T=106210 14010 0 0 $X=106070 $Y=13300
X187 6 VIA1_C_CDNS_724652923740 $T=106210 38730 0 0 $X=106070 $Y=38020
X188 3 VIA2_C_CDNS_724652923741 $T=7870 104220 0 0 $X=6900 $Y=103560
X189 3 VIA2_C_CDNS_724652923741 $T=7870 131040 0 0 $X=6900 $Y=130380
X190 6 VIA2_C_CDNS_724652923741 $T=11050 15465 0 0 $X=10080 $Y=14805
X191 6 VIA2_C_CDNS_724652923741 $T=11050 40105 0 0 $X=10080 $Y=39445
X192 6 VIA2_C_CDNS_724652923741 $T=29650 15465 0 0 $X=28680 $Y=14805
X193 6 VIA2_C_CDNS_724652923741 $T=29650 40105 0 0 $X=28680 $Y=39445
X194 14 VIA2_C_CDNS_724652923741 $T=38035 56445 0 0 $X=37065 $Y=55785
X195 14 VIA2_C_CDNS_724652923741 $T=38035 89245 0 0 $X=37065 $Y=88585
X196 12 VIA2_C_CDNS_724652923741 $T=40315 58225 0 0 $X=39345 $Y=57565
X197 12 VIA2_C_CDNS_724652923741 $T=40315 85685 0 0 $X=39345 $Y=85025
X198 14 VIA2_C_CDNS_724652923741 $T=40420 12230 0 0 $X=39450 $Y=11570
X199 14 VIA2_C_CDNS_724652923741 $T=40420 42290 0 0 $X=39450 $Y=41630
X200 6 VIA2_C_CDNS_724652923741 $T=42700 14010 0 0 $X=41730 $Y=13350
X201 6 VIA2_C_CDNS_724652923741 $T=42700 38730 0 0 $X=41730 $Y=38070
X202 3 VIA2_C_CDNS_724652923741 $T=43570 104220 0 0 $X=42600 $Y=103560
X203 3 VIA2_C_CDNS_724652923741 $T=43570 131040 0 0 $X=42600 $Y=130380
X204 12 VIA2_C_CDNS_724652923741 $T=107055 58225 0 0 $X=106085 $Y=57565
X205 12 VIA2_C_CDNS_724652923741 $T=107055 85685 0 0 $X=106085 $Y=85025
X206 6 VIA2_C_CDNS_724652923741 $T=108020 14010 0 0 $X=107050 $Y=13350
X207 6 VIA2_C_CDNS_724652923741 $T=108020 38730 0 0 $X=107050 $Y=38070
X208 13 VIA2_C_CDNS_724652923741 $T=109335 54665 0 0 $X=108365 $Y=54005
X209 13 VIA2_C_CDNS_724652923741 $T=109335 87465 0 0 $X=108365 $Y=86805
X210 13 VIA2_C_CDNS_724652923741 $T=110300 10450 0 0 $X=109330 $Y=9790
X211 13 VIA2_C_CDNS_724652923741 $T=110300 40510 0 0 $X=109330 $Y=39850
X212 4 VIA1_C_CDNS_724652923742 $T=10135 89745 0 0 $X=9995 $Y=89555
X213 5 VIA1_C_CDNS_724652923742 $T=10845 66505 0 0 $X=10705 $Y=66315
X214 4 VIA1_C_CDNS_724652923742 $T=11675 89745 0 0 $X=11535 $Y=89555
X215 5 VIA1_C_CDNS_724652923742 $T=12385 66505 0 0 $X=12245 $Y=66315
X216 4 VIA1_C_CDNS_724652923742 $T=13215 89745 0 0 $X=13075 $Y=89555
X217 5 VIA1_C_CDNS_724652923742 $T=13925 66505 0 0 $X=13785 $Y=66315
X218 4 VIA1_C_CDNS_724652923742 $T=14755 89745 0 0 $X=14615 $Y=89555
X219 5 VIA1_C_CDNS_724652923742 $T=15465 66505 0 0 $X=15325 $Y=66315
X220 2 VIA1_C_CDNS_724652923742 $T=15870 27855 0 0 $X=15730 $Y=27665
X221 2 VIA1_C_CDNS_724652923742 $T=18110 27855 0 0 $X=17970 $Y=27665
X222 2 VIA1_C_CDNS_724652923742 $T=20350 27855 0 0 $X=20210 $Y=27665
X223 2 VIA1_C_CDNS_724652923742 $T=22590 27855 0 0 $X=22450 $Y=27665
X224 5 VIA1_C_CDNS_724652923742 $T=23230 66505 0 0 $X=23090 $Y=66315
X225 5 VIA1_C_CDNS_724652923742 $T=24770 66505 0 0 $X=24630 $Y=66315
X226 2 VIA1_C_CDNS_724652923742 $T=24830 27855 0 0 $X=24690 $Y=27665
X227 5 VIA1_C_CDNS_724652923742 $T=26310 66505 0 0 $X=26170 $Y=66315
X228 5 VIA1_C_CDNS_724652923742 $T=27850 66505 0 0 $X=27710 $Y=66315
X229 1 VIA2_C_CDNS_724652923743 $T=5840 100660 0 0 $X=5130 $Y=100000
X230 1 VIA2_C_CDNS_724652923743 $T=5840 134600 0 0 $X=5130 $Y=133940
X231 2 VIA2_C_CDNS_724652923743 $T=7240 13685 0 0 $X=6530 $Y=13025
X232 2 VIA2_C_CDNS_724652923743 $T=7240 43665 0 0 $X=6530 $Y=43005
X233 8 VIA2_C_CDNS_724652923743 $T=9020 11905 0 0 $X=8310 $Y=11245
X234 8 VIA2_C_CDNS_724652923743 $T=9020 41885 0 0 $X=8310 $Y=41225
X235 11 VIA2_C_CDNS_724652923743 $T=31680 45445 0 0 $X=30970 $Y=44785
X236 10 VIA2_C_CDNS_724652923743 $T=33460 10125 0 0 $X=32750 $Y=9465
X237 9 VIA2_C_CDNS_724652923743 $T=45600 102440 0 0 $X=44890 $Y=101780
X238 9 VIA2_C_CDNS_724652923743 $T=45600 136380 0 0 $X=44890 $Y=135720
X239 7 VIA2_C_CDNS_724652923743 $T=47380 98880 0 0 $X=46670 $Y=98220
X240 7 VIA2_C_CDNS_724652923743 $T=47380 132820 0 0 $X=46670 $Y=132160
X241 1 VIA2_C_CDNS_724652923744 $T=5840 117700 0 0 $X=5130 $Y=117560
X242 2 VIA2_C_CDNS_724652923744 $T=7240 27855 0 0 $X=6530 $Y=27715
X243 1 VIA1_C_CDNS_724652923745 $T=13400 117700 0 0 $X=13000 $Y=117510
X244 1 VIA1_C_CDNS_724652923745 $T=15640 117700 0 0 $X=15240 $Y=117510
X245 1 VIA1_C_CDNS_724652923745 $T=17880 117700 0 0 $X=17480 $Y=117510
X246 1 VIA1_C_CDNS_724652923745 $T=20120 117700 0 0 $X=19720 $Y=117510
X247 1 VIA1_C_CDNS_724652923745 $T=22360 117700 0 0 $X=21960 $Y=117510
X248 4 VIA1_C_CDNS_724652923745 $T=23940 89745 0 0 $X=23540 $Y=89555
X249 1 VIA1_C_CDNS_724652923745 $T=24600 117700 0 0 $X=24200 $Y=117510
X250 4 VIA1_C_CDNS_724652923745 $T=25480 89745 0 0 $X=25080 $Y=89555
X251 1 VIA1_C_CDNS_724652923745 $T=26840 117700 0 0 $X=26440 $Y=117510
X252 4 VIA1_C_CDNS_724652923745 $T=27020 89745 0 0 $X=26620 $Y=89555
X253 4 VIA1_C_CDNS_724652923745 $T=28560 89745 0 0 $X=28160 $Y=89555
X254 1 VIA1_C_CDNS_724652923745 $T=29080 117700 0 0 $X=28680 $Y=117510
X255 1 VIA1_C_CDNS_724652923745 $T=31320 117700 0 0 $X=30920 $Y=117510
X256 1 VIA1_C_CDNS_724652923745 $T=33560 117700 0 0 $X=33160 $Y=117510
X257 1 VIA1_C_CDNS_724652923745 $T=35800 117700 0 0 $X=35400 $Y=117510
X258 1 VIA1_C_CDNS_724652923745 $T=38040 117700 0 0 $X=37640 $Y=117510
X259 17 VIA1_C_CDNS_724652923745 $T=51305 71565 0 0 $X=50905 $Y=71375
X260 18 VIA1_C_CDNS_724652923745 $T=52955 72345 0 0 $X=52555 $Y=72155
X261 14 VIA1_C_CDNS_724652923745 $T=53520 26400 0 0 $X=53120 $Y=26210
X262 17 VIA1_C_CDNS_724652923745 $T=58085 71565 0 0 $X=57685 $Y=71375
X263 18 VIA1_C_CDNS_724652923745 $T=58765 72345 0 0 $X=58365 $Y=72155
X264 14 VIA1_C_CDNS_724652923745 $T=59760 26400 0 0 $X=59360 $Y=26210
X265 19 VIA1_C_CDNS_724652923745 $T=62155 117840 0 0 $X=61755 $Y=117650
X266 17 VIA1_C_CDNS_724652923745 $T=63785 71565 0 0 $X=63385 $Y=71375
X267 18 VIA1_C_CDNS_724652923745 $T=65435 72345 0 0 $X=65035 $Y=72155
X268 14 VIA1_C_CDNS_724652923745 $T=66000 26400 0 0 $X=65600 $Y=26210
X269 19 VIA1_C_CDNS_724652923745 $T=68395 117840 0 0 $X=67995 $Y=117650
X270 17 VIA1_C_CDNS_724652923745 $T=70565 71565 0 0 $X=70165 $Y=71375
X271 18 VIA1_C_CDNS_724652923745 $T=71245 72345 0 0 $X=70845 $Y=72155
X272 14 VIA1_C_CDNS_724652923745 $T=72240 26400 0 0 $X=71840 $Y=26210
X273 17 VIA1_C_CDNS_724652923745 $T=76265 71565 0 0 $X=75865 $Y=71375
X274 18 VIA1_C_CDNS_724652923745 $T=77915 72345 0 0 $X=77515 $Y=72155
X275 14 VIA1_C_CDNS_724652923745 $T=78480 26400 0 0 $X=78080 $Y=26210
X276 15 VIA1_C_CDNS_724652923745 $T=81575 136880 0 0 $X=81175 $Y=136690
X277 17 VIA1_C_CDNS_724652923745 $T=83045 71565 0 0 $X=82645 $Y=71375
X278 18 VIA1_C_CDNS_724652923745 $T=83725 72345 0 0 $X=83325 $Y=72155
X279 14 VIA1_C_CDNS_724652923745 $T=84720 26400 0 0 $X=84320 $Y=26210
X280 15 VIA1_C_CDNS_724652923745 $T=87815 136880 0 0 $X=87415 $Y=136690
X281 17 VIA1_C_CDNS_724652923745 $T=88745 71565 0 0 $X=88345 $Y=71375
X282 18 VIA1_C_CDNS_724652923745 $T=90395 72345 0 0 $X=89995 $Y=72155
X283 14 VIA1_C_CDNS_724652923745 $T=90960 26400 0 0 $X=90560 $Y=26210
X284 17 VIA1_C_CDNS_724652923745 $T=95525 71565 0 0 $X=95125 $Y=71375
X285 18 VIA1_C_CDNS_724652923745 $T=96205 72345 0 0 $X=95805 $Y=72155
X286 13 VIA1_C_CDNS_724652923745 $T=96290 114275 0 0 $X=95890 $Y=114085
X287 14 VIA1_C_CDNS_724652923745 $T=97200 26400 0 0 $X=96800 $Y=26210
X288 13 VIA1_C_CDNS_724652923745 $T=97830 114275 0 0 $X=97430 $Y=114085
X289 7 VIA1_C_CDNS_724652923745 $T=98460 136920 0 0 $X=98060 $Y=136730
X290 13 VIA1_C_CDNS_724652923745 $T=99370 114275 0 0 $X=98970 $Y=114085
X291 20 VIA1_C_CDNS_724652923745 $T=100700 136140 0 0 $X=100300 $Y=135950
X292 13 VIA1_C_CDNS_724652923745 $T=100910 114275 0 0 $X=100510 $Y=114085
X293 3 VIA1_C_CDNS_724652923746 $T=59385 131570 0 0 $X=59245 $Y=130600
X294 19 VIA1_C_CDNS_724652923746 $T=64925 133850 0 0 $X=64785 $Y=132880
X295 3 VIA1_C_CDNS_724652923746 $T=65625 131570 0 0 $X=65485 $Y=130600
X296 18 VIA1_C_CDNS_724652923746 $T=71165 136130 0 0 $X=71025 $Y=135160
X297 10 VIA1_C_CDNS_724652923746 $T=97690 123640 0 0 $X=97550 $Y=122670
X298 15 VIA1_C_CDNS_724652923746 $T=99230 121360 0 0 $X=99090 $Y=120390
X299 10 VIA1_C_CDNS_724652923746 $T=99930 123640 0 0 $X=99790 $Y=122670
X300 16 VIA1_C_CDNS_724652923746 $T=101470 119080 0 0 $X=101330 $Y=118110
X301 6 VIA1_C_CDNS_724652923748 $T=95520 101635 0 0 $X=95120 $Y=100665
X302 7 VIA1_C_CDNS_724652923748 $T=97060 99355 0 0 $X=96660 $Y=98385
X303 6 VIA1_C_CDNS_724652923748 $T=98600 101635 0 0 $X=98200 $Y=100665
X304 7 VIA1_C_CDNS_724652923748 $T=100140 99355 0 0 $X=99740 $Y=98385
X305 6 VIA1_C_CDNS_724652923748 $T=101680 101635 0 0 $X=101280 $Y=100665
X306 6 VIA2_C_CDNS_724652923749 $T=20350 6575 0 0 $X=16220 $Y=5565
X307 6 VIA2_C_CDNS_724652923749 $T=75360 6055 0 0 $X=71230 $Y=5045
X308 6 VIA1_C_CDNS_7246529237410 $T=20350 6575 0 0 $X=16220 $Y=5565
X309 6 VIA1_C_CDNS_7246529237410 $T=75360 6055 0 0 $X=71230 $Y=5045
X310 3 VIA1_C_CDNS_7246529237412 $T=6000 138620 0 0 $X=4210 $Y=137870
X311 3 VIA1_C_CDNS_7246529237412 $T=47220 138620 0 0 $X=45430 $Y=137870
X312 3 VIA1_C_CDNS_7246529237412 $T=59055 138620 0 0 $X=57265 $Y=137870
X313 3 VIA1_C_CDNS_7246529237412 $T=84905 138620 0 0 $X=83115 $Y=137870
X314 3 VIA1_C_CDNS_7246529237414 $T=110725 50485 0 0 $X=110235 $Y=47655
X315 3 VIA1_C_CDNS_7246529237414 $T=119195 38515 0 0 $X=118705 $Y=35685
X316 7 VIA1_C_CDNS_7246529237415 $T=118805 88080 0 0 $X=118315 $Y=86030
X317 7 VIA1_C_CDNS_7246529237415 $T=118805 136570 0 0 $X=118315 $Y=134520
X318 17 VIA1_C_CDNS_7246529237415 $T=208665 49725 0 0 $X=208175 $Y=47675
X319 18 VIA1_C_CDNS_7246529237415 $T=208725 98250 0 0 $X=208235 $Y=96200
X320 1 VIA2_C_CDNS_7246529237420 $T=9255 74485 0 0 $X=8505 $Y=73735
X321 8 VIA2_C_CDNS_7246529237420 $T=22885 54255 0 0 $X=22135 $Y=53505
X322 21 VIA1_C_CDNS_7246529237422 $T=296735 11275 0 0 $X=296245 $Y=7145
X323 17 VIA1_C_CDNS_7246529237422 $T=296735 36110 0 0 $X=296245 $Y=31980
X324 21 VIA1_C_CDNS_7246529237424 $T=307595 14520 0 0 $X=307405 $Y=10480
X325 21 VIA1_C_CDNS_7246529237424 $T=307595 31270 0 0 $X=307405 $Y=27230
X326 21 VIA1_C_CDNS_7246529237424 $T=307595 48020 0 0 $X=307405 $Y=43980
X327 21 VIA1_C_CDNS_7246529237424 $T=307595 64770 0 0 $X=307405 $Y=60730
X328 21 VIA1_C_CDNS_7246529237424 $T=307595 81520 0 0 $X=307405 $Y=77480
X329 21 VIA1_C_CDNS_7246529237424 $T=307595 98270 0 0 $X=307405 $Y=94230
X330 21 VIA1_C_CDNS_7246529237424 $T=307595 115020 0 0 $X=307405 $Y=110980
X331 21 VIA1_C_CDNS_7246529237424 $T=307595 131770 0 0 $X=307405 $Y=127730
X332 21 VIA1_C_CDNS_7246529237424 $T=324350 14520 0 0 $X=324160 $Y=10480
X333 21 VIA1_C_CDNS_7246529237424 $T=324350 31270 0 0 $X=324160 $Y=27230
X334 21 VIA1_C_CDNS_7246529237424 $T=324350 48020 0 0 $X=324160 $Y=43980
X335 21 VIA1_C_CDNS_7246529237424 $T=324350 81520 0 0 $X=324160 $Y=77480
X336 21 VIA1_C_CDNS_7246529237424 $T=324350 98270 0 0 $X=324160 $Y=94230
X337 21 VIA1_C_CDNS_7246529237424 $T=324350 115020 0 0 $X=324160 $Y=110980
X338 21 VIA1_C_CDNS_7246529237424 $T=324350 131770 0 0 $X=324160 $Y=127730
X339 21 VIA1_C_CDNS_7246529237424 $T=341105 14520 0 0 $X=340915 $Y=10480
X340 21 VIA1_C_CDNS_7246529237424 $T=341105 31270 0 0 $X=340915 $Y=27230
X341 21 VIA1_C_CDNS_7246529237424 $T=341105 48020 0 0 $X=340915 $Y=43980
X342 21 VIA1_C_CDNS_7246529237424 $T=341105 64770 0 0 $X=340915 $Y=60730
X343 21 VIA1_C_CDNS_7246529237424 $T=341105 81520 0 0 $X=340915 $Y=77480
X344 21 VIA1_C_CDNS_7246529237424 $T=341105 98270 0 0 $X=340915 $Y=94230
X345 21 VIA1_C_CDNS_7246529237424 $T=341105 115020 0 0 $X=340915 $Y=110980
X346 21 VIA1_C_CDNS_7246529237424 $T=341105 131770 0 0 $X=340915 $Y=127730
X347 21 VIA1_C_CDNS_7246529237424 $T=357860 14520 0 0 $X=357670 $Y=10480
X348 21 VIA1_C_CDNS_7246529237424 $T=357860 31270 0 0 $X=357670 $Y=27230
X349 21 VIA1_C_CDNS_7246529237424 $T=357860 48020 0 0 $X=357670 $Y=43980
X350 21 VIA1_C_CDNS_7246529237424 $T=357860 64770 0 0 $X=357670 $Y=60730
X351 21 VIA1_C_CDNS_7246529237424 $T=357860 81520 0 0 $X=357670 $Y=77480
X352 21 VIA1_C_CDNS_7246529237424 $T=357860 98270 0 0 $X=357670 $Y=94230
X353 21 VIA1_C_CDNS_7246529237424 $T=357860 115020 0 0 $X=357670 $Y=110980
X354 21 VIA1_C_CDNS_7246529237424 $T=357860 131770 0 0 $X=357670 $Y=127730
X355 7 VIA2_C_CDNS_7246529237429 $T=118800 136695 0 0 $X=118310 $Y=134645
X356 18 VIA2_C_CDNS_7246529237429 $T=208725 98250 0 0 $X=208235 $Y=96200
X357 1 4 4 3 6 pe3_CDNS_724652923740 $T=9635 78185 0 0 $X=8125 $Y=77155
X358 9 4 12 3 6 pe3_CDNS_724652923740 $T=23440 78185 0 0 $X=21930 $Y=77155
X359 2 5 5 6 ne3_CDNS_724652923741 $T=10345 55405 0 0 $X=9545 $Y=55005
X360 8 5 4 6 ne3_CDNS_724652923741 $T=22730 55545 0 0 $X=21930 $Y=55145
X361 6 13 7 6 ne3_CDNS_724652923741 $T=95790 103175 0 0 $X=94990 $Y=102775
X362 17 21 6 rpp1k1_3_CDNS_724652923742 $T=287735 7255 1 180 $X=159445 $Y=7035
X363 7 22 6 rpp1k1_3_CDNS_724652923743 $T=123895 47740 0 0 $X=118735 $Y=47520
X364 6 6 6 6 ne3_CDNS_724652923744 $T=13130 16755 0 0 $X=12330 $Y=16355
X365 6 6 6 6 ne3_CDNS_724652923744 $T=13130 38815 1 0 $X=12330 $Y=28245
X366 6 2 8 6 ne3_CDNS_724652923744 $T=15370 16755 0 0 $X=14570 $Y=16355
X367 6 2 2 6 ne3_CDNS_724652923744 $T=15370 38815 1 0 $X=14570 $Y=28245
X368 6 2 2 6 ne3_CDNS_724652923744 $T=17610 16755 0 0 $X=16810 $Y=16355
X369 6 2 8 6 ne3_CDNS_724652923744 $T=17610 38815 1 0 $X=16810 $Y=28245
X370 6 2 10 6 ne3_CDNS_724652923744 $T=19850 16755 0 0 $X=19050 $Y=16355
X371 6 2 11 6 ne3_CDNS_724652923744 $T=19850 38815 1 0 $X=19050 $Y=28245
X372 6 2 8 6 ne3_CDNS_724652923744 $T=22090 16755 0 0 $X=21290 $Y=16355
X373 6 2 2 6 ne3_CDNS_724652923744 $T=22090 38815 1 0 $X=21290 $Y=28245
X374 6 2 2 6 ne3_CDNS_724652923744 $T=24330 16755 0 0 $X=23530 $Y=16355
X375 6 2 8 6 ne3_CDNS_724652923744 $T=24330 38815 1 0 $X=23530 $Y=28245
X376 6 6 6 6 ne3_CDNS_724652923744 $T=26570 16755 0 0 $X=25770 $Y=16355
X377 6 6 6 6 ne3_CDNS_724652923744 $T=26570 38815 1 0 $X=25770 $Y=28245
X378 10 7 15 6 ne3_CDNS_724652923744 $T=97960 125180 0 0 $X=97160 $Y=124780
X379 10 20 16 6 ne3_CDNS_724652923744 $T=100200 125180 0 0 $X=99400 $Y=124780
X380 12 12 12 3 6 pe3_CDNS_724652923746 $T=43105 60145 0 0 $X=41595 $Y=59115
X381 12 12 12 3 6 pe3_CDNS_724652923746 $T=43105 83765 1 0 $X=41595 $Y=72735
X382 12 18 13 3 6 pe3_CDNS_724652923746 $T=49345 60145 0 0 $X=47835 $Y=59115
X383 12 17 14 3 6 pe3_CDNS_724652923746 $T=49345 83765 1 0 $X=47835 $Y=72735
X384 12 17 14 3 6 pe3_CDNS_724652923746 $T=55585 60145 0 0 $X=54075 $Y=59115
X385 12 18 13 3 6 pe3_CDNS_724652923746 $T=55585 83765 1 0 $X=54075 $Y=72735
X386 3 19 19 3 6 pe3_CDNS_724652923746 $T=59655 129400 1 0 $X=58145 $Y=118370
X387 12 18 13 3 6 pe3_CDNS_724652923746 $T=61825 60145 0 0 $X=60315 $Y=59115
X388 12 17 14 3 6 pe3_CDNS_724652923746 $T=61825 83765 1 0 $X=60315 $Y=72735
X389 3 19 18 3 6 pe3_CDNS_724652923746 $T=65895 129400 1 0 $X=64385 $Y=118370
X390 12 17 14 3 6 pe3_CDNS_724652923746 $T=68065 60145 0 0 $X=66555 $Y=59115
X391 12 18 13 3 6 pe3_CDNS_724652923746 $T=68065 83765 1 0 $X=66555 $Y=72735
X392 12 18 13 3 6 pe3_CDNS_724652923746 $T=74305 60145 0 0 $X=72795 $Y=59115
X393 12 17 14 3 6 pe3_CDNS_724652923746 $T=74305 83765 1 0 $X=72795 $Y=72735
X394 3 15 15 3 6 pe3_CDNS_724652923746 $T=79075 125320 0 0 $X=77565 $Y=124290
X395 12 17 14 3 6 pe3_CDNS_724652923746 $T=80545 60145 0 0 $X=79035 $Y=59115
X396 12 18 13 3 6 pe3_CDNS_724652923746 $T=80545 83765 1 0 $X=79035 $Y=72735
X397 3 15 16 3 6 pe3_CDNS_724652923746 $T=85315 125320 0 0 $X=83805 $Y=124290
X398 12 18 13 3 6 pe3_CDNS_724652923746 $T=86785 60145 0 0 $X=85275 $Y=59115
X399 12 17 14 3 6 pe3_CDNS_724652923746 $T=86785 83765 1 0 $X=85275 $Y=72735
X400 12 17 14 3 6 pe3_CDNS_724652923746 $T=93025 60145 0 0 $X=91515 $Y=59115
X401 12 18 13 3 6 pe3_CDNS_724652923746 $T=93025 83765 1 0 $X=91515 $Y=72735
X402 12 12 12 3 6 pe3_CDNS_724652923746 $T=99265 60145 0 0 $X=97755 $Y=59115
X403 12 12 12 3 6 pe3_CDNS_724652923746 $T=99265 83765 1 0 $X=97755 $Y=72735
X404 19 16 11 3 6 pe3_CDNS_724652923747 $T=62750 104210 0 0 $X=61240 $Y=103180
X405 6 20 6 ne3_CDNS_724652923748 $T=110195 126990 0 0 $X=109395 $Y=126590
X406 20 23 6 ne3_CDNS_724652923748 $T=110195 130510 0 0 $X=109395 $Y=130110
X407 23 3 6 ne3_CDNS_724652923748 $T=110195 134045 0 0 $X=109395 $Y=133645
X408 3 3 3 6 pe3_CDNS_724652923749 $T=10660 106140 0 0 $X=9150 $Y=105110
X409 3 3 3 6 pe3_CDNS_724652923749 $T=10660 129120 1 0 $X=9150 $Y=118090
X410 3 1 7 6 pe3_CDNS_724652923749 $T=12900 106140 0 0 $X=11390 $Y=105110
X411 3 1 7 6 pe3_CDNS_724652923749 $T=12900 129120 1 0 $X=11390 $Y=118090
X412 3 1 7 6 pe3_CDNS_724652923749 $T=15140 106140 0 0 $X=13630 $Y=105110
X413 3 1 7 6 pe3_CDNS_724652923749 $T=15140 129120 1 0 $X=13630 $Y=118090
X414 3 1 9 6 pe3_CDNS_724652923749 $T=17380 106140 0 0 $X=15870 $Y=105110
X415 3 1 1 6 pe3_CDNS_724652923749 $T=17380 129120 1 0 $X=15870 $Y=118090
X416 3 1 7 6 pe3_CDNS_724652923749 $T=19620 106140 0 0 $X=18110 $Y=105110
X417 3 1 7 6 pe3_CDNS_724652923749 $T=19620 129120 1 0 $X=18110 $Y=118090
X418 3 1 7 6 pe3_CDNS_724652923749 $T=21860 106140 0 0 $X=20350 $Y=105110
X419 3 1 7 6 pe3_CDNS_724652923749 $T=21860 129120 1 0 $X=20350 $Y=118090
X420 3 1 1 6 pe3_CDNS_724652923749 $T=24100 106140 0 0 $X=22590 $Y=105110
X421 3 1 9 6 pe3_CDNS_724652923749 $T=24100 129120 1 0 $X=22590 $Y=118090
X422 3 1 9 6 pe3_CDNS_724652923749 $T=26340 106140 0 0 $X=24830 $Y=105110
X423 3 1 1 6 pe3_CDNS_724652923749 $T=26340 129120 1 0 $X=24830 $Y=118090
X424 3 1 7 6 pe3_CDNS_724652923749 $T=28580 106140 0 0 $X=27070 $Y=105110
X425 3 1 7 6 pe3_CDNS_724652923749 $T=28580 129120 1 0 $X=27070 $Y=118090
X426 3 1 7 6 pe3_CDNS_724652923749 $T=30820 106140 0 0 $X=29310 $Y=105110
X427 3 1 7 6 pe3_CDNS_724652923749 $T=30820 129120 1 0 $X=29310 $Y=118090
X428 3 1 1 6 pe3_CDNS_724652923749 $T=33060 106140 0 0 $X=31550 $Y=105110
X429 3 1 9 6 pe3_CDNS_724652923749 $T=33060 129120 1 0 $X=31550 $Y=118090
X430 3 1 7 6 pe3_CDNS_724652923749 $T=35300 106140 0 0 $X=33790 $Y=105110
X431 3 1 7 6 pe3_CDNS_724652923749 $T=35300 129120 1 0 $X=33790 $Y=118090
X432 3 1 7 6 pe3_CDNS_724652923749 $T=37540 106140 0 0 $X=36030 $Y=105110
X433 3 1 7 6 pe3_CDNS_724652923749 $T=37540 129120 1 0 $X=36030 $Y=118090
X434 3 3 3 6 pe3_CDNS_724652923749 $T=39780 106140 0 0 $X=38270 $Y=105110
X435 3 3 3 6 pe3_CDNS_724652923749 $T=39780 129120 1 0 $X=38270 $Y=118090
X436 6 6 6 ne3_CDNS_7246529237410 $T=44780 15300 0 0 $X=43980 $Y=14900
X437 6 6 6 ne3_CDNS_7246529237410 $T=44780 37440 1 0 $X=43980 $Y=26870
X438 6 14 14 ne3_CDNS_7246529237410 $T=51020 15300 0 0 $X=50220 $Y=14900
X439 6 14 13 ne3_CDNS_7246529237410 $T=51020 37440 1 0 $X=50220 $Y=26870
X440 6 14 13 ne3_CDNS_7246529237410 $T=57260 15300 0 0 $X=56460 $Y=14900
X441 6 14 14 ne3_CDNS_7246529237410 $T=57260 37440 1 0 $X=56460 $Y=26870
X442 6 14 14 ne3_CDNS_7246529237410 $T=63500 15300 0 0 $X=62700 $Y=14900
X443 6 14 13 ne3_CDNS_7246529237410 $T=63500 37440 1 0 $X=62700 $Y=26870
X444 6 14 13 ne3_CDNS_7246529237410 $T=69740 15300 0 0 $X=68940 $Y=14900
X445 6 14 14 ne3_CDNS_7246529237410 $T=69740 37440 1 0 $X=68940 $Y=26870
X446 6 14 14 ne3_CDNS_7246529237410 $T=75980 15300 0 0 $X=75180 $Y=14900
X447 6 14 13 ne3_CDNS_7246529237410 $T=75980 37440 1 0 $X=75180 $Y=26870
X448 6 14 13 ne3_CDNS_7246529237410 $T=82220 15300 0 0 $X=81420 $Y=14900
X449 6 14 14 ne3_CDNS_7246529237410 $T=82220 37440 1 0 $X=81420 $Y=26870
X450 6 14 14 ne3_CDNS_7246529237410 $T=88460 15300 0 0 $X=87660 $Y=14900
X451 6 14 13 ne3_CDNS_7246529237410 $T=88460 37440 1 0 $X=87660 $Y=26870
X452 6 14 13 ne3_CDNS_7246529237410 $T=94700 15300 0 0 $X=93900 $Y=14900
X453 6 14 14 ne3_CDNS_7246529237410 $T=94700 37440 1 0 $X=93900 $Y=26870
X454 6 6 6 ne3_CDNS_7246529237410 $T=100940 15300 0 0 $X=100140 $Y=14900
X455 6 6 6 ne3_CDNS_7246529237410 $T=100940 37440 1 0 $X=100140 $Y=26870
X456 7 24 6 rpp1k1_3_CDNS_7246529237411 $T=123895 96235 0 0 $X=118735 $Y=96015
X457 22 17 6 rpp1k1_3_CDNS_7246529237411 $T=213685 47740 0 0 $X=208525 $Y=47520
X458 24 18 6 rpp1k1_3_CDNS_7246529237411 $T=213685 96235 0 0 $X=208525 $Y=96015
Q0 6 6 21 qpvc3 $X=302595 $Y=9520 $dt=2
Q1 6 6 21 qpvc3 $X=302595 $Y=26270 $dt=2
Q2 6 6 21 qpvc3 $X=302595 $Y=43020 $dt=2
Q3 6 6 21 qpvc3 $X=302595 $Y=59770 $dt=2
Q4 6 6 21 qpvc3 $X=302595 $Y=76520 $dt=2
Q5 6 6 21 qpvc3 $X=302595 $Y=93270 $dt=2
Q6 6 6 21 qpvc3 $X=302595 $Y=110020 $dt=2
Q7 6 6 21 qpvc3 $X=302595 $Y=126770 $dt=2
Q8 6 6 21 qpvc3 $X=319350 $Y=9520 $dt=2
Q9 6 6 21 qpvc3 $X=319350 $Y=26270 $dt=2
Q10 6 6 21 qpvc3 $X=319350 $Y=43020 $dt=2
Q11 6 6 18 qpvc3 $X=319350 $Y=59770 $dt=2
Q12 6 6 21 qpvc3 $X=319350 $Y=76520 $dt=2
Q13 6 6 21 qpvc3 $X=319350 $Y=93270 $dt=2
Q14 6 6 21 qpvc3 $X=319350 $Y=110020 $dt=2
Q15 6 6 21 qpvc3 $X=319350 $Y=126770 $dt=2
Q16 6 6 21 qpvc3 $X=336105 $Y=9520 $dt=2
Q17 6 6 21 qpvc3 $X=336105 $Y=26270 $dt=2
Q18 6 6 21 qpvc3 $X=336105 $Y=43020 $dt=2
Q19 6 6 21 qpvc3 $X=336105 $Y=59770 $dt=2
Q20 6 6 21 qpvc3 $X=336105 $Y=76520 $dt=2
Q21 6 6 21 qpvc3 $X=336105 $Y=93270 $dt=2
Q22 6 6 21 qpvc3 $X=336105 $Y=110020 $dt=2
Q23 6 6 21 qpvc3 $X=336105 $Y=126770 $dt=2
Q24 6 6 21 qpvc3 $X=352860 $Y=9520 $dt=2
Q25 6 6 21 qpvc3 $X=352860 $Y=26270 $dt=2
Q26 6 6 21 qpvc3 $X=352860 $Y=43020 $dt=2
Q27 6 6 21 qpvc3 $X=352860 $Y=59770 $dt=2
Q28 6 6 21 qpvc3 $X=352860 $Y=76520 $dt=2
Q29 6 6 21 qpvc3 $X=352860 $Y=93270 $dt=2
Q30 6 6 21 qpvc3 $X=352860 $Y=110020 $dt=2
Q31 6 6 21 qpvc3 $X=352860 $Y=126770 $dt=2
D32 6 3 p_dnw AREA=1.07147e-09 PJ=0.0001732 perimeter=0.0001732 $X=3950 $Y=96990 $dt=3
D33 6 3 p_dnw AREA=2.50005e-10 PJ=8.653e-05 perimeter=8.653e-05 $X=6985 $Y=72595 $dt=3
D34 6 3 p_dnw AREA=1.35123e-09 PJ=0.00022788 perimeter=0.00022788 $X=35895 $Y=52775 $dt=3
D35 6 3 p_dnw AREA=3.30547e-10 PJ=0.00010554 perimeter=0.00010554 $X=57005 $Y=102040 $dt=3
D36 6 3 p_dnw AREA=1.64117e-10 PJ=7.372e-05 perimeter=7.372e-05 $X=76425 $Y=117950 $dt=3
D37 6 3 p_dnw AREA=1.17512e-09 PJ=0.00013712 perimeter=0.00013712 $X=119255 $Y=7325 $dt=3
D38 6 3 p_dnw3 AREA=3.99668e-10 PJ=0 perimeter=0 $X=9150 $Y=105110 $dt=4
D39 6 3 p_dnw3 AREA=3.99668e-10 PJ=0 perimeter=0 $X=9150 $Y=118090 $dt=4
D40 6 3 p_dnw3 AREA=7.74011e-10 PJ=0 perimeter=0 $X=41595 $Y=59115 $dt=4
D41 6 3 p_dnw3 AREA=7.74011e-10 PJ=0 perimeter=0 $X=41595 $Y=72735 $dt=4
D42 6 3 p_dnw3 AREA=1.71976e-10 PJ=0 perimeter=0 $X=58145 $Y=118370 $dt=4
D43 6 3 p_dnw3 AREA=1.71976e-10 PJ=0 perimeter=0 $X=77565 $Y=124290 $dt=4
C44 13 7 area=9e-10 perimeter=0.00012 $[cmm5t] $X=121395 $Y=9465 $dt=6
.ends bandgap_su
