* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : emir_test_1                                  *
* Netlisted  : Wed Jul 17 08:24:21 2024                     *
* PVS Version: 23.10-p043 Mon Oct 2 18:09:08 PDT 2023      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 R(rpp1k1) rpp1k1_2 p1trm(POS) p1trm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_CDNS_721219056720                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_CDNS_721219056720 2 3
** N=3 EP=2 FDC=1
R0 2 3 L=2.5e-05 W=5e-06 $[rpp1k1] $X=0 $Y=0 $dt=0
.ends rpp1k1_CDNS_721219056720

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: emir_test_1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt emir_test_1 gnda vdda
** N=3 EP=2 FDC=3
X0 gnda vdda rpp1k1_CDNS_721219056720 $T=314165 13865 0 180 $X=288225 $Y=8645
X1 gnda vdda rpp1k1_CDNS_721219056720 $T=314165 23360 0 180 $X=288225 $Y=18140
X2 gnda vdda rpp1k1_CDNS_721219056720 $T=314165 34615 0 180 $X=288225 $Y=29395
.ends emir_test_1
