* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : bandgap_su                                   *
* Netlisted  : Mon Aug 26 08:15:29 2024                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(ne3) nem ndiff(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 1 MP(pe3) pem pdiff(D) p1trm(G) pdiff(S) nwtrm(B)
*.DEVTMPLT 2 Q(qpvc3) qpvmc bulk(C) nwtrm(B) pdiff(E)
*.DEVTMPLT 3 D(p_dnw) p_dnw bulk(POS) nwtrm(NEG)
*.DEVTMPLT 4 D(p_dnw3) p_dnwm bulk(POS) nwtrm(NEG)
*.DEVTMPLT 5 R(rpp1k1_3) rpp1k1_s p1trm(POS) p1trm(NEG) bulk(SUB)
*.DEVTMPLT 6 C(cmm5t) cmim capm(POS) m4trm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724652923740                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724652923740 1 2 3 4 5
** N=5 EP=5 FDC=5
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=1
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=1
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=1
D4 5 4 p_dnw3 AREA=1.04198e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=4
.ends pe3_CDNS_724652923740

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724652923741                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724652923741 1 2 3 4
** N=4 EP=4 FDC=4
M0 3 2 1 4 ne3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
M1 1 2 3 4 ne3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=0
M2 3 2 1 4 ne3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=0
M3 1 2 3 4 ne3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=0
.ends ne3_CDNS_724652923741

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_724652923742                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_724652923742 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.0005215 W=8e-06 $[rpp1k1_3] $SUB=3 $X=-8220 $Y=0 $dt=5
.ends rpp1k1_3_CDNS_724652923742

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_724652923743                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_724652923743 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.00082283 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=5
.ends rpp1k1_3_CDNS_724652923743

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724652923744                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724652923744 1 2 3 4
** N=4 EP=4 FDC=1
M0 3 2 1 4 ne3 L=1e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
.ends ne3_CDNS_724652923744

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724652923746                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724652923746 1 2 3 4
*.DEVICECLIMB
** N=5 EP=4 FDC=1
M0 3 2 1 4 pe3 L=5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_724652923746

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724652923747                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724652923747 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 3 2 1 4 pe3 L=5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
D1 5 4 p_dnw3 AREA=9.67212e-11 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=4
.ends pe3_CDNS_724652923747

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724652923748                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724652923748 1 2 3
** N=3 EP=3 FDC=1
M0 2 2 1 3 ne3 L=2e-06 W=1e-06 AD=4.8e-13 AS=4.8e-13 PD=2.96e-06 PS=2.96e-06 $X=0 $Y=0 $dt=0
.ends ne3_CDNS_724652923748

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724652923749                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724652923749 1 2 3
*.DEVICECLIMB
** N=4 EP=3 FDC=1
M0 3 2 1 1 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_724652923749

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7246529237410                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7246529237410 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
.ends ne3_CDNS_7246529237410

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7246529237411                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7246529237411 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.00082283 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=5
.ends rpp1k1_3_CDNS_7246529237411

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: bandgap_su                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt bandgap_su BIAS GNDA OUT VDD3A
** N=24 EP=4 FDC=165
X357 1 4 4 VDD3A GNDA pe3_CDNS_724652923740 $T=9635 78185 0 0 $X=8125 $Y=77155
X358 9 4 12 VDD3A GNDA pe3_CDNS_724652923740 $T=23440 78185 0 0 $X=21930 $Y=77155
X359 2 BIAS BIAS GNDA ne3_CDNS_724652923741 $T=10345 55405 0 0 $X=9545 $Y=55005
X360 8 BIAS 4 GNDA ne3_CDNS_724652923741 $T=22730 55545 0 0 $X=21930 $Y=55145
X361 GNDA 13 OUT GNDA ne3_CDNS_724652923741 $T=95790 103175 0 0 $X=94990 $Y=102775
X362 17 21 GNDA rpp1k1_3_CDNS_724652923742 $T=287735 7255 1 180 $X=159445 $Y=7035
X363 OUT 22 GNDA rpp1k1_3_CDNS_724652923743 $T=123895 47740 0 0 $X=118735 $Y=47520
X364 GNDA GNDA GNDA GNDA ne3_CDNS_724652923744 $T=13130 16755 0 0 $X=12330 $Y=16355
X365 GNDA GNDA GNDA GNDA ne3_CDNS_724652923744 $T=13130 38815 1 0 $X=12330 $Y=28245
X366 GNDA 2 8 GNDA ne3_CDNS_724652923744 $T=15370 16755 0 0 $X=14570 $Y=16355
X367 GNDA 2 2 GNDA ne3_CDNS_724652923744 $T=15370 38815 1 0 $X=14570 $Y=28245
X368 GNDA 2 2 GNDA ne3_CDNS_724652923744 $T=17610 16755 0 0 $X=16810 $Y=16355
X369 GNDA 2 8 GNDA ne3_CDNS_724652923744 $T=17610 38815 1 0 $X=16810 $Y=28245
X370 GNDA 2 10 GNDA ne3_CDNS_724652923744 $T=19850 16755 0 0 $X=19050 $Y=16355
X371 GNDA 2 11 GNDA ne3_CDNS_724652923744 $T=19850 38815 1 0 $X=19050 $Y=28245
X372 GNDA 2 8 GNDA ne3_CDNS_724652923744 $T=22090 16755 0 0 $X=21290 $Y=16355
X373 GNDA 2 2 GNDA ne3_CDNS_724652923744 $T=22090 38815 1 0 $X=21290 $Y=28245
X374 GNDA 2 2 GNDA ne3_CDNS_724652923744 $T=24330 16755 0 0 $X=23530 $Y=16355
X375 GNDA 2 8 GNDA ne3_CDNS_724652923744 $T=24330 38815 1 0 $X=23530 $Y=28245
X376 GNDA GNDA GNDA GNDA ne3_CDNS_724652923744 $T=26570 16755 0 0 $X=25770 $Y=16355
X377 GNDA GNDA GNDA GNDA ne3_CDNS_724652923744 $T=26570 38815 1 0 $X=25770 $Y=28245
X378 10 OUT 15 GNDA ne3_CDNS_724652923744 $T=97960 125180 0 0 $X=97160 $Y=124780
X379 10 20 16 GNDA ne3_CDNS_724652923744 $T=100200 125180 0 0 $X=99400 $Y=124780
X380 12 12 12 VDD3A pe3_CDNS_724652923746 $T=43105 60145 0 0 $X=41595 $Y=59115
X381 12 12 12 VDD3A pe3_CDNS_724652923746 $T=43105 83765 1 0 $X=41595 $Y=72735
X382 12 18 13 VDD3A pe3_CDNS_724652923746 $T=49345 60145 0 0 $X=47835 $Y=59115
X383 12 17 14 VDD3A pe3_CDNS_724652923746 $T=49345 83765 1 0 $X=47835 $Y=72735
X384 12 17 14 VDD3A pe3_CDNS_724652923746 $T=55585 60145 0 0 $X=54075 $Y=59115
X385 12 18 13 VDD3A pe3_CDNS_724652923746 $T=55585 83765 1 0 $X=54075 $Y=72735
X386 VDD3A 19 19 VDD3A pe3_CDNS_724652923746 $T=59655 129400 1 0 $X=58145 $Y=118370
X387 12 18 13 VDD3A pe3_CDNS_724652923746 $T=61825 60145 0 0 $X=60315 $Y=59115
X388 12 17 14 VDD3A pe3_CDNS_724652923746 $T=61825 83765 1 0 $X=60315 $Y=72735
X389 VDD3A 19 18 VDD3A pe3_CDNS_724652923746 $T=65895 129400 1 0 $X=64385 $Y=118370
X390 12 17 14 VDD3A pe3_CDNS_724652923746 $T=68065 60145 0 0 $X=66555 $Y=59115
X391 12 18 13 VDD3A pe3_CDNS_724652923746 $T=68065 83765 1 0 $X=66555 $Y=72735
X392 12 18 13 VDD3A pe3_CDNS_724652923746 $T=74305 60145 0 0 $X=72795 $Y=59115
X393 12 17 14 VDD3A pe3_CDNS_724652923746 $T=74305 83765 1 0 $X=72795 $Y=72735
X394 VDD3A 15 15 VDD3A pe3_CDNS_724652923746 $T=79075 125320 0 0 $X=77565 $Y=124290
X395 12 17 14 VDD3A pe3_CDNS_724652923746 $T=80545 60145 0 0 $X=79035 $Y=59115
X396 12 18 13 VDD3A pe3_CDNS_724652923746 $T=80545 83765 1 0 $X=79035 $Y=72735
X397 VDD3A 15 16 VDD3A pe3_CDNS_724652923746 $T=85315 125320 0 0 $X=83805 $Y=124290
X398 12 18 13 VDD3A pe3_CDNS_724652923746 $T=86785 60145 0 0 $X=85275 $Y=59115
X399 12 17 14 VDD3A pe3_CDNS_724652923746 $T=86785 83765 1 0 $X=85275 $Y=72735
X400 12 17 14 VDD3A pe3_CDNS_724652923746 $T=93025 60145 0 0 $X=91515 $Y=59115
X401 12 18 13 VDD3A pe3_CDNS_724652923746 $T=93025 83765 1 0 $X=91515 $Y=72735
X402 12 12 12 VDD3A pe3_CDNS_724652923746 $T=99265 60145 0 0 $X=97755 $Y=59115
X403 12 12 12 VDD3A pe3_CDNS_724652923746 $T=99265 83765 1 0 $X=97755 $Y=72735
X404 19 16 11 VDD3A GNDA pe3_CDNS_724652923747 $T=62750 104210 0 0 $X=61240 $Y=103180
X405 GNDA 20 GNDA ne3_CDNS_724652923748 $T=110195 126990 0 0 $X=109395 $Y=126590
X406 20 23 GNDA ne3_CDNS_724652923748 $T=110195 130510 0 0 $X=109395 $Y=130110
X407 23 VDD3A GNDA ne3_CDNS_724652923748 $T=110195 134045 0 0 $X=109395 $Y=133645
X408 VDD3A VDD3A VDD3A pe3_CDNS_724652923749 $T=10660 106140 0 0 $X=9150 $Y=105110
X409 VDD3A VDD3A VDD3A pe3_CDNS_724652923749 $T=10660 129120 1 0 $X=9150 $Y=118090
X410 VDD3A 1 OUT pe3_CDNS_724652923749 $T=12900 106140 0 0 $X=11390 $Y=105110
X411 VDD3A 1 OUT pe3_CDNS_724652923749 $T=12900 129120 1 0 $X=11390 $Y=118090
X412 VDD3A 1 OUT pe3_CDNS_724652923749 $T=15140 106140 0 0 $X=13630 $Y=105110
X413 VDD3A 1 OUT pe3_CDNS_724652923749 $T=15140 129120 1 0 $X=13630 $Y=118090
X414 VDD3A 1 9 pe3_CDNS_724652923749 $T=17380 106140 0 0 $X=15870 $Y=105110
X415 VDD3A 1 1 pe3_CDNS_724652923749 $T=17380 129120 1 0 $X=15870 $Y=118090
X416 VDD3A 1 OUT pe3_CDNS_724652923749 $T=19620 106140 0 0 $X=18110 $Y=105110
X417 VDD3A 1 OUT pe3_CDNS_724652923749 $T=19620 129120 1 0 $X=18110 $Y=118090
X418 VDD3A 1 OUT pe3_CDNS_724652923749 $T=21860 106140 0 0 $X=20350 $Y=105110
X419 VDD3A 1 OUT pe3_CDNS_724652923749 $T=21860 129120 1 0 $X=20350 $Y=118090
X420 VDD3A 1 1 pe3_CDNS_724652923749 $T=24100 106140 0 0 $X=22590 $Y=105110
X421 VDD3A 1 9 pe3_CDNS_724652923749 $T=24100 129120 1 0 $X=22590 $Y=118090
X422 VDD3A 1 9 pe3_CDNS_724652923749 $T=26340 106140 0 0 $X=24830 $Y=105110
X423 VDD3A 1 1 pe3_CDNS_724652923749 $T=26340 129120 1 0 $X=24830 $Y=118090
X424 VDD3A 1 OUT pe3_CDNS_724652923749 $T=28580 106140 0 0 $X=27070 $Y=105110
X425 VDD3A 1 OUT pe3_CDNS_724652923749 $T=28580 129120 1 0 $X=27070 $Y=118090
X426 VDD3A 1 OUT pe3_CDNS_724652923749 $T=30820 106140 0 0 $X=29310 $Y=105110
X427 VDD3A 1 OUT pe3_CDNS_724652923749 $T=30820 129120 1 0 $X=29310 $Y=118090
X428 VDD3A 1 1 pe3_CDNS_724652923749 $T=33060 106140 0 0 $X=31550 $Y=105110
X429 VDD3A 1 9 pe3_CDNS_724652923749 $T=33060 129120 1 0 $X=31550 $Y=118090
X430 VDD3A 1 OUT pe3_CDNS_724652923749 $T=35300 106140 0 0 $X=33790 $Y=105110
X431 VDD3A 1 OUT pe3_CDNS_724652923749 $T=35300 129120 1 0 $X=33790 $Y=118090
X432 VDD3A 1 OUT pe3_CDNS_724652923749 $T=37540 106140 0 0 $X=36030 $Y=105110
X433 VDD3A 1 OUT pe3_CDNS_724652923749 $T=37540 129120 1 0 $X=36030 $Y=118090
X434 VDD3A VDD3A VDD3A pe3_CDNS_724652923749 $T=39780 106140 0 0 $X=38270 $Y=105110
X435 VDD3A VDD3A VDD3A pe3_CDNS_724652923749 $T=39780 129120 1 0 $X=38270 $Y=118090
X436 GNDA GNDA GNDA ne3_CDNS_7246529237410 $T=44780 15300 0 0 $X=43980 $Y=14900
X437 GNDA GNDA GNDA ne3_CDNS_7246529237410 $T=44780 37440 1 0 $X=43980 $Y=26870
X438 GNDA 14 14 ne3_CDNS_7246529237410 $T=51020 15300 0 0 $X=50220 $Y=14900
X439 GNDA 14 13 ne3_CDNS_7246529237410 $T=51020 37440 1 0 $X=50220 $Y=26870
X440 GNDA 14 13 ne3_CDNS_7246529237410 $T=57260 15300 0 0 $X=56460 $Y=14900
X441 GNDA 14 14 ne3_CDNS_7246529237410 $T=57260 37440 1 0 $X=56460 $Y=26870
X442 GNDA 14 14 ne3_CDNS_7246529237410 $T=63500 15300 0 0 $X=62700 $Y=14900
X443 GNDA 14 13 ne3_CDNS_7246529237410 $T=63500 37440 1 0 $X=62700 $Y=26870
X444 GNDA 14 13 ne3_CDNS_7246529237410 $T=69740 15300 0 0 $X=68940 $Y=14900
X445 GNDA 14 14 ne3_CDNS_7246529237410 $T=69740 37440 1 0 $X=68940 $Y=26870
X446 GNDA 14 14 ne3_CDNS_7246529237410 $T=75980 15300 0 0 $X=75180 $Y=14900
X447 GNDA 14 13 ne3_CDNS_7246529237410 $T=75980 37440 1 0 $X=75180 $Y=26870
X448 GNDA 14 13 ne3_CDNS_7246529237410 $T=82220 15300 0 0 $X=81420 $Y=14900
X449 GNDA 14 14 ne3_CDNS_7246529237410 $T=82220 37440 1 0 $X=81420 $Y=26870
X450 GNDA 14 14 ne3_CDNS_7246529237410 $T=88460 15300 0 0 $X=87660 $Y=14900
X451 GNDA 14 13 ne3_CDNS_7246529237410 $T=88460 37440 1 0 $X=87660 $Y=26870
X452 GNDA 14 13 ne3_CDNS_7246529237410 $T=94700 15300 0 0 $X=93900 $Y=14900
X453 GNDA 14 14 ne3_CDNS_7246529237410 $T=94700 37440 1 0 $X=93900 $Y=26870
X454 GNDA GNDA GNDA ne3_CDNS_7246529237410 $T=100940 15300 0 0 $X=100140 $Y=14900
X455 GNDA GNDA GNDA ne3_CDNS_7246529237410 $T=100940 37440 1 0 $X=100140 $Y=26870
X456 OUT 24 GNDA rpp1k1_3_CDNS_7246529237411 $T=123895 96235 0 0 $X=118735 $Y=96015
X457 22 17 GNDA rpp1k1_3_CDNS_7246529237411 $T=213685 47740 0 0 $X=208525 $Y=47520
X458 24 18 GNDA rpp1k1_3_CDNS_7246529237411 $T=213685 96235 0 0 $X=208525 $Y=96015
Q0 GNDA GNDA 21 qpvc3 $X=302595 $Y=9520 $dt=2
Q1 GNDA GNDA 21 qpvc3 $X=302595 $Y=26270 $dt=2
Q2 GNDA GNDA 21 qpvc3 $X=302595 $Y=43020 $dt=2
Q3 GNDA GNDA 21 qpvc3 $X=302595 $Y=59770 $dt=2
Q4 GNDA GNDA 21 qpvc3 $X=302595 $Y=76520 $dt=2
Q5 GNDA GNDA 21 qpvc3 $X=302595 $Y=93270 $dt=2
Q6 GNDA GNDA 21 qpvc3 $X=302595 $Y=110020 $dt=2
Q7 GNDA GNDA 21 qpvc3 $X=302595 $Y=126770 $dt=2
Q8 GNDA GNDA 21 qpvc3 $X=319350 $Y=9520 $dt=2
Q9 GNDA GNDA 21 qpvc3 $X=319350 $Y=26270 $dt=2
Q10 GNDA GNDA 21 qpvc3 $X=319350 $Y=43020 $dt=2
Q11 GNDA GNDA 18 qpvc3 $X=319350 $Y=59770 $dt=2
Q12 GNDA GNDA 21 qpvc3 $X=319350 $Y=76520 $dt=2
Q13 GNDA GNDA 21 qpvc3 $X=319350 $Y=93270 $dt=2
Q14 GNDA GNDA 21 qpvc3 $X=319350 $Y=110020 $dt=2
Q15 GNDA GNDA 21 qpvc3 $X=319350 $Y=126770 $dt=2
Q16 GNDA GNDA 21 qpvc3 $X=336105 $Y=9520 $dt=2
Q17 GNDA GNDA 21 qpvc3 $X=336105 $Y=26270 $dt=2
Q18 GNDA GNDA 21 qpvc3 $X=336105 $Y=43020 $dt=2
Q19 GNDA GNDA 21 qpvc3 $X=336105 $Y=59770 $dt=2
Q20 GNDA GNDA 21 qpvc3 $X=336105 $Y=76520 $dt=2
Q21 GNDA GNDA 21 qpvc3 $X=336105 $Y=93270 $dt=2
Q22 GNDA GNDA 21 qpvc3 $X=336105 $Y=110020 $dt=2
Q23 GNDA GNDA 21 qpvc3 $X=336105 $Y=126770 $dt=2
Q24 GNDA GNDA 21 qpvc3 $X=352860 $Y=9520 $dt=2
Q25 GNDA GNDA 21 qpvc3 $X=352860 $Y=26270 $dt=2
Q26 GNDA GNDA 21 qpvc3 $X=352860 $Y=43020 $dt=2
Q27 GNDA GNDA 21 qpvc3 $X=352860 $Y=59770 $dt=2
Q28 GNDA GNDA 21 qpvc3 $X=352860 $Y=76520 $dt=2
Q29 GNDA GNDA 21 qpvc3 $X=352860 $Y=93270 $dt=2
Q30 GNDA GNDA 21 qpvc3 $X=352860 $Y=110020 $dt=2
Q31 GNDA GNDA 21 qpvc3 $X=352860 $Y=126770 $dt=2
D32 GNDA VDD3A p_dnw AREA=1.07147e-09 PJ=0.0001732 perimeter=0.0001732 $X=3950 $Y=96990 $dt=3
D33 GNDA VDD3A p_dnw AREA=2.50005e-10 PJ=8.653e-05 perimeter=8.653e-05 $X=6985 $Y=72595 $dt=3
D34 GNDA VDD3A p_dnw AREA=1.35123e-09 PJ=0.00022788 perimeter=0.00022788 $X=35895 $Y=52775 $dt=3
D35 GNDA VDD3A p_dnw AREA=3.30547e-10 PJ=0.00010554 perimeter=0.00010554 $X=57005 $Y=102040 $dt=3
D36 GNDA VDD3A p_dnw AREA=1.64117e-10 PJ=7.372e-05 perimeter=7.372e-05 $X=76425 $Y=117950 $dt=3
D37 GNDA VDD3A p_dnw AREA=1.17512e-09 PJ=0.00013712 perimeter=0.00013712 $X=119255 $Y=7325 $dt=3
D38 GNDA VDD3A p_dnw3 AREA=3.99668e-10 PJ=0 perimeter=0 $X=9150 $Y=105110 $dt=4
D39 GNDA VDD3A p_dnw3 AREA=3.99668e-10 PJ=0 perimeter=0 $X=9150 $Y=118090 $dt=4
D40 GNDA VDD3A p_dnw3 AREA=7.74011e-10 PJ=0 perimeter=0 $X=41595 $Y=59115 $dt=4
D41 GNDA VDD3A p_dnw3 AREA=7.74011e-10 PJ=0 perimeter=0 $X=41595 $Y=72735 $dt=4
D42 GNDA VDD3A p_dnw3 AREA=1.71976e-10 PJ=0 perimeter=0 $X=58145 $Y=118370 $dt=4
D43 GNDA VDD3A p_dnw3 AREA=1.71976e-10 PJ=0 perimeter=0 $X=77565 $Y=124290 $dt=4
C44 13 OUT area=9e-10 perimeter=0.00012 $[cmm5t] $X=121395 $Y=9465 $dt=6
.ends bandgap_su
