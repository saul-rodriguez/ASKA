* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : emir_test_2                                  *
* Netlisted  : Wed Aug  7 04:01:24 2024                     *
* PVS Version: 23.10-p043 Mon Oct 2 18:09:08 PDT 2023      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 R(rpp1k1) rpp1k1_2 p1trm(POS) p1trm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_723017679630                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_723017679630 1 2
** N=2 EP=2 FDC=0
.ends VIATP_C_CDNS_723017679630

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_723017679631                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_723017679631 1 2
** N=2 EP=2 FDC=0
.ends VIA3_C_CDNS_723017679631

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_723017679632                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_723017679632 1 2
** N=2 EP=2 FDC=0
.ends VIA2_C_CDNS_723017679632

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_723017679633                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_723017679633 1 2
** N=2 EP=2 FDC=0
.ends VIA1_C_CDNS_723017679633

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_CDNS_723017679630                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_CDNS_723017679630 1 2 3
** N=3 EP=3 FDC=1
R0 2 3 L=2.5e-05 W=5e-06 $[rpp1k1] $X=0 $Y=0 $dt=0
.ends rpp1k1_CDNS_723017679630

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: emir_test_2                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt emir_test_2 3 2
** N=4 EP=2 FDC=7
X0 1 2 VIATP_C_CDNS_723017679630 $T=2825 71645 0 0 $X=2090 $Y=53870
X1 1 2 VIATP_C_CDNS_723017679630 $T=289560 71645 0 0 $X=288825 $Y=53870
X2 1 2 VIA3_C_CDNS_723017679631 $T=2825 71645 0 0 $X=2090 $Y=53770
X3 1 2 VIA3_C_CDNS_723017679631 $T=289560 71645 0 0 $X=288825 $Y=53770
X4 1 2 VIA2_C_CDNS_723017679632 $T=2825 71645 0 0 $X=2290 $Y=53970
X5 1 2 VIA2_C_CDNS_723017679632 $T=289560 71645 0 0 $X=289025 $Y=53970
X6 1 2 VIA1_C_CDNS_723017679633 $T=2825 71645 0 0 $X=2290 $Y=53970
X7 1 2 VIA1_C_CDNS_723017679633 $T=289560 71645 0 0 $X=289025 $Y=53970
X8 1 3 2 rpp1k1_CDNS_723017679630 $T=314165 13865 0 180 $X=288225 $Y=8645
X9 1 3 2 rpp1k1_CDNS_723017679630 $T=314165 23360 0 180 $X=288225 $Y=18140
X10 1 3 2 rpp1k1_CDNS_723017679630 $T=314165 34615 0 180 $X=288225 $Y=29395
X11 1 2 3 rpp1k1_CDNS_723017679630 $T=290815 57190 0 0 $X=289875 $Y=56970
X12 1 2 3 rpp1k1_CDNS_723017679630 $T=290815 65265 0 0 $X=289875 $Y=65045
X13 1 2 3 rpp1k1_CDNS_723017679630 $T=290815 72930 0 0 $X=289875 $Y=72710
X14 1 2 3 rpp1k1_CDNS_723017679630 $T=290815 80325 0 0 $X=289875 $Y=80105
.ends emir_test_2
