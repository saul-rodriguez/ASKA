************************************************************************
* auCdl Netlist:
* 
* Library Name:  ASKA_BANDGAP
* Top Cell Name: bandgap_su
* View Name:     schematic
* Netlisted on:  Aug 26 08:15:24 2024
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.LDD
*.SCALE METER
.PARAM



************************************************************************
* Library Name: ASKA_BANDGAP
* Cell Name:    bandgap_su
* View Name:    schematic
************************************************************************

.SUBCKT bandgap_su BIAS GNDA OUT VDD3A
*.PININFO BIAS:B GNDA:B OUT:B VDD3A:B
MM29 GNDA GNDA GNDA GNDA NE3 W=10u L=5u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM25 net21 net21 GNDA GNDA NE3 W=1u L=2u M=1.0 AD=4.8e-13 AS=4.8e-13 
+ PD=2.96e-06 PS=2.96e-06 NRD=0.27 NRS=0.27
MM24 VDD3A VDD3A net22 GNDA NE3 W=1u L=2u M=1.0 AD=4.8e-13 AS=4.8e-13 
+ PD=2.96e-06 PS=2.96e-06 NRD=0.27 NRS=0.27
MM23 net22 net22 net21 GNDA NE3 W=1u L=2u M=1.0 AD=4.8e-13 AS=4.8e-13 
+ PD=2.96e-06 PS=2.96e-06 NRD=0.27 NRS=0.27
MM26 GNDA GNDA GNDA GNDA NE3 W=10u L=1u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM17 net12 net21 net7 GNDA NE3 W=10u L=1u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM16 net10 OUT net7 GNDA NE3 W=10u L=1u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM15 net7 net6 GNDA GNDA NE3 W=10u L=1u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM14 net1 net6 GNDA GNDA NE3 W=10u L=1u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM13 OUT net17 GNDA GNDA NE3 W=10u L=1u M=4.0 AD=2.7e-12 AS=3.75e-12 
+ PD=1.054e-05 PS=1.575e-05 NRD=0.027 NRS=0.027
MM11 net3 BIAS net2 GNDA NE3 W=10u L=1u M=4.0 AD=2.7e-12 AS=3.75e-12 
+ PD=1.054e-05 PS=1.575e-05 NRD=0.027 NRS=0.027
MM9 BIAS BIAS net6 GNDA NE3 W=10u L=1u M=4.0 AD=2.7e-12 AS=3.75e-12 
+ PD=1.054e-05 PS=1.575e-05 NRD=0.027 NRS=0.027
MM8 net2 net6 GNDA GNDA NE3 W=10u L=1u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM7 net6 net6 GNDA GNDA NE3 W=10u L=1u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM4 net15 net15 GNDA GNDA NE3 W=10u L=5u M=8.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM2 net17 net15 GNDA GNDA NE3 W=10u L=5u M=8.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM28 A A A VDD3A PE3 W=10u L=5u M=4.0 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 
+ PS=2.096e-05 NRD=0.027 NRS=0.027
MM27 VDD3A VDD3A VDD3A VDD3A PE3 W=10u L=1u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM22 net11 net20 VDD3A VDD3A PE3 W=10u L=5u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM21 net1 net12 net20 VDD3A PE3 W=10u L=5u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM20 net20 net20 VDD3A VDD3A PE3 W=10u L=5u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM19 net12 net10 VDD3A VDD3A PE3 W=10u L=5u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM18 net10 net10 VDD3A VDD3A PE3 W=10u L=5u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM12 OUT net16 VDD3A VDD3A PE3 W=10u L=1u M=16.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM6 net3 net3 net16 VDD3A PE3 W=10u L=1u M=4.0 AD=2.7e-12 AS=3.75e-12 
+ PD=1.054e-05 PS=1.575e-05 NRD=0.027 NRS=0.027
MM1 A net3 net14 VDD3A PE3 W=10u L=1u M=4.0 AD=2.7e-12 AS=3.75e-12 
+ PD=1.054e-05 PS=1.575e-05 NRD=0.027 NRS=0.027
MM0 net16 net16 VDD3A VDD3A PE3 W=10u L=1u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM10 net14 net16 VDD3A VDD3A PE3 W=10u L=1u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM5 net17 net11 A VDD3A PE3 W=10u L=5u M=8.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM3 net15 net23 A VDD3A PE3 W=10u L=5u M=8.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
QQ6 GNDA GNDA net11 QPVC3 1e-10 M=1
QQ5 GNDA GNDA net9 QPVC3 1e-10 M=31
RR11 net5 OUT 200.032K $SUB=GNDA $[RPP1K1_3] $W=4u $L=822.83u M=1
RR10 net8 OUT 200.032K $SUB=GNDA $[RPP1K1_3] $W=4u $L=822.83u M=1
RR8 net23 net5 200.032K $SUB=GNDA $[RPP1K1_3] $W=4u $L=822.83u M=1
RR7 net9 net23 63000 $SUB=GNDA $[RPP1K1_3] $W=8u $L=521.5u M=1
RR6 net11 net8 200.032K $SUB=GNDA $[RPP1K1_3] $W=4u $L=822.83u M=1
CC1 net17 OUT $[CMM5T] area=9e-10 perimeter=120.00000u M=1
.ENDS

