* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : del_test                                     *
* Netlisted  : Fri Aug 23 11:27:24 2024                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(ne3) nem ndiff(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 1 MP(pe3) pem pdiff(D) p1trm(G) pdiff(S) nwtrm(B)
*.DEVTMPLT 2 D(p_dnw3) p_dnwm bulk(POS) nwtrm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724405238730                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724405238730 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724405238730

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_724405238731                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_724405238731 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_724405238731

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_724405238732                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_724405238732 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_724405238732

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: IN_3VX2                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt IN_3VX2 1 2 3 4
** N=4 EP=4 FDC=5
M0 4 3 2 2 ne3 L=3.5e-07 W=4.8e-07 AD=1.296e-13 AS=4.408e-13 PD=1.02e-06 PS=3.52e-06 $X=500 $Y=1070 $dt=0
M1 2 3 4 2 ne3 L=3.5e-07 W=4.8e-07 AD=4.408e-13 AS=1.296e-13 PD=3.52e-06 PS=1.02e-06 $X=1390 $Y=1070 $dt=0
M2 4 3 1 1 pe3 L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=8.151e-13 PD=1.87971e-06 PS=4.50971e-06 $X=560 $Y=2410 $dt=1
M3 1 3 4 1 pe3 L=3.00472e-07 W=1.45971e-06 AD=8.01e-13 AS=2.751e-13 PD=4.48971e-06 PS=1.87971e-06 $X=1400 $Y=2410 $dt=1
D4 2 1 p_dnw3 AREA=9.734e-12 PJ=1.248e-05 perimeter=1.248e-05 $X=-430 $Y=1980 $dt=2
.ends IN_3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: IN_3VX4                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt IN_3VX4 1 2 3 4
** N=4 EP=4 FDC=8
M0 2 4 3 2 ne3 L=3.5e-07 W=8e-07 AD=4.148e-13 AS=3.84e-13 PD=1.98e-06 PS=2.56e-06 $X=620 $Y=750 $dt=0
M1 3 4 2 2 ne3 L=3.5e-07 W=8e-07 AD=2.16e-13 AS=4.148e-13 PD=1.34e-06 PS=1.98e-06 $X=1710 $Y=750 $dt=0
M2 2 4 3 2 ne3 L=3.5e-07 W=8e-07 AD=9.852e-13 AS=2.16e-13 PD=4.14e-06 PS=1.34e-06 $X=2600 $Y=750 $dt=0
M3 3 4 1 1 pe3 L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=5.79287e-13 PD=1.86506e-06 PS=3.69506e-06 $X=475 $Y=2410 $dt=1
M4 1 4 3 1 pe3 L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=1315 $Y=2410 $dt=1
M5 3 4 1 1 pe3 L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=1865 $Y=2410 $dt=1
M6 1 4 3 1 pe3 L=3.00566e-07 W=1.47006e-06 AD=1.48669e-12 AS=2.54913e-13 PD=5.27506e-06 PS=1.86506e-06 $X=2705 $Y=2410 $dt=1
D7 2 1 p_dnw3 AREA=1.50092e-11 PJ=1.584e-05 perimeter=1.584e-05 $X=-430 $Y=1980 $dt=2
.ends IN_3VX4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: del_test                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt del_test 3 7 5 6 2
** N=7 EP=5 FDC=26
X0 1 VIA1_C_CDNS_724405238730 $T=-930 64845 0 0 $X=-1120 $Y=64705
X1 1 VIA1_C_CDNS_724405238730 $T=2998795 64845 0 0 $X=2998605 $Y=64705
X2 1 VIA2_C_CDNS_724405238731 $T=-60 64845 0 0 $X=-250 $Y=64705
X3 1 VIA2_C_CDNS_724405238731 $T=2997705 64845 0 0 $X=2997515 $Y=64705
X4 1 VIA3_C_CDNS_724405238732 $T=755 64845 0 0 $X=565 $Y=64705
X5 1 VIA3_C_CDNS_724405238732 $T=2996520 64845 0 0 $X=2996330 $Y=64705
X6 2 3 4 5 IN_3VX2 $T=2999540 25295 0 0 $X=2999110 $Y=24655
X7 2 3 1 6 IN_3VX2 $T=2999540 66790 1 0 $X=2999110 $Y=61670
X8 2 3 4 7 IN_3VX4 $T=-4380 25295 0 0 $X=-4810 $Y=24655
X9 2 3 1 7 IN_3VX4 $T=-4380 66790 1 0 $X=-4810 $Y=61670
.ends del_test
