* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : ne3i_test3                                   *
* Netlisted  : Sun Jun 23 12:47:38 2024                     *
* PVS Version: 23.10-p043 Mon Oct 2 18:09:08 PDT 2023      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 NE3I_6() nemi_6 ndiff(D) p1trm(G) ndiff(S) pwitrm(B) dnwtrm(NW) bulk(SB)
*.DEVTMPLT 1 D(p_ddnw) p_ddnw bulk(POS) dnwtrm(NEG)
*.DEVTMPLT 2 D(p_dipdnwmv) p_dipwmv pwitrm(POS) dnwtrm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NE3I_6                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NE3I_6 D G S B NW SB
.ends NE3I_6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3i_6_CDNS_719161253260                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3i_6_CDNS_719161253260 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=1
X0 1 2 3 1 4 5 NE3I_6 w=1e-05 l=2e-06 as=4.8e-12 ad=4.8e-12 ps=2.096e-05 pd=2.096e-05 $X=0 $Y=0 $dt=0
.ends ne3i_6_CDNS_719161253260

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3i_test3                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3i_test3 GNDA INN INP OU1 OU2 VDDA
** N=7 EP=6 FDC=6
X20 1 INN OU2 VDDA GNDA ne3i_6_CDNS_719161253260 $T=12675 18045 0 0 $X=8615 $Y=13595
X21 1 INP OU1 VDDA GNDA ne3i_6_CDNS_719161253260 $T=12675 42845 1 0 $X=8615 $Y=28275
X22 1 INP OU1 VDDA GNDA ne3i_6_CDNS_719161253260 $T=16075 18045 0 0 $X=12015 $Y=13595
X23 1 INN OU2 VDDA GNDA ne3i_6_CDNS_719161253260 $T=16075 42845 1 0 $X=12015 $Y=28275
D0 GNDA VDDA p_ddnw AREA=5.02014e-10 PJ=0.0001046 perimeter=0.0001046 $X=7345 $Y=12325 $dt=1
D1 1 VDDA p_dipdnwmv AREA=1.58594e-10 PJ=7.38e-05 perimeter=7.38e-05 $X=11195 $Y=16175 $dt=2
.ends ne3i_test3
