************************************************************************
* auCdl Netlist:
* 
* Library Name:  ASKA_BIAS
* Top Cell Name: bias
* View Name:     schematic
* Netlisted on:  Aug 26 08:36:55 2024
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.LDD
*.SCALE METER
.PARAM



************************************************************************
* Library Name: ASKA_CONSTANT_GM
* Cell Name:    constant_gm
* View Name:    schematic
************************************************************************

.SUBCKT constant_gm GNDA OUT1 OUT2 OUT3 VDD3
*.PININFO GNDA:B OUT1:B OUT2:B OUT3:B VDD3:B
MM1 net1 net1 net13 GNDA NE3 W=10u L=2.5u M=2.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM0 net24 net1 net23 GNDA NE3 W=10u L=2.5u M=2.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM17 VDD3 VDD3 VDD3 VDD3 PE3 W=10u L=2.5u M=5.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM16 net47 net17 VDD3 VDD3 PE3 W=10u L=2.5u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM15 OUT3 net24 net47 VDD3 PE3 W=10u L=2.5u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM14 net2 net2 net24 net24 PE3 W=2u L=10u M=1.0 AD=9.6e-13 AS=9.6e-13 
+ PD=4.96e-06 PS=4.96e-06 NRD=0.135 NRS=0.135
MM13 net40 net17 VDD3 VDD3 PE3 W=10u L=2.5u M=2.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM11 OUT2 net24 net40 VDD3 PE3 W=10u L=2.5u M=2.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM8 net1 net1 net2 net2 PE3 W=2u L=10u M=1.0 AD=9.6e-13 AS=9.6e-13 PD=4.96e-06 
+ PS=4.96e-06 NRD=0.135 NRS=0.135
MM7 OUT1 net24 net30 VDD3 PE3 W=10u L=2.5u M=2.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM6 net30 net17 VDD3 VDD3 PE3 W=10u L=2.5u M=2.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM5 net1 net24 net18 VDD3 PE3 W=10u L=2.5u M=2.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM3 net24 net24 net17 VDD3 PE3 W=10u L=2.5u M=2.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM9 net18 net17 VDD3 VDD3 PE3 W=10u L=2.5u M=2.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM12 net17 net17 VDD3 VDD3 PE3 W=10u L=2.5u M=2.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
RR3 GNDA net25 69999.7 $SUB=VDD3 $[RPP1K1_3] $W=4u $L=287.8u M=1
XM4 net13 net13 GNDA GNDA VDD3 GNDA / ne3i_6 W=10u L=2.5u M=2.0 AD=2.7e-12 
+ AS=4.8e-12 NRD=0.027 NRS=0.027 PD=1.054e-05 PS=2.096e-05 par1=2.0
XM2 net23 net13 net25 net25 VDD3 GNDA / ne3i_6 W=10u L=2.5u M=8.0 AD=2.7e-12 
+ AS=3.225e-12 NRD=0.027 NRS=0.027 PD=1.054e-05 PS=1.3145e-05 par1=8.0
.ENDS

************************************************************************
* Library Name: ASKA_REF_BIAS
* Cell Name:    ref_bias
* View Name:    schematic
************************************************************************

.SUBCKT ref_bias BIAS GNDA OUT1 OUT2 RES_BIAS VDDA VREF
*.PININFO BIAS:B GNDA:B OUT1:B OUT2:B RES_BIAS:B VDDA:B VREF:B
XM7 COM COM COM COM VDDA GNDA / ne3i_6 W=10u L=2u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ NRD=0.027 NRS=0.027 PD=2.096e-05 PS=2.096e-05 par1=4.0
XM12 net4 VREF COM COM VDDA GNDA / ne3i_6 W=10u L=2u M=14.0 AD=4.8e-12 
+ AS=4.8e-12 NRD=0.027 NRS=0.027 PD=2.096e-05 PS=2.096e-05 par1=14.0
XM24 net6 RES_BIAS COM COM VDDA GNDA / ne3i_6 W=10u L=2u M=14.0 AD=4.8e-12 
+ AS=4.8e-12 NRD=0.027 NRS=0.027 PD=2.096e-05 PS=2.096e-05 par1=14.0
MM10 GNDA GNDA GNDA GNDA NE3 W=10u L=5u M=5.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM9 BIAS BIAS net123 GNDA NE3 W=10u L=2u M=8.0 AD=2.7e-12 AS=3.225e-12 
+ PD=1.054e-05 PS=1.3145e-05 NRD=0.027 NRS=0.027
MM8 COM BIAS net5 GNDA NE3 W=10u L=2u M=8.0 AD=2.7e-12 AS=3.225e-12 
+ PD=1.054e-05 PS=1.3145e-05 NRD=0.027 NRS=0.027
MM26 net7 net123 GNDA GNDA NE3 W=10u L=5u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM13 net123 net123 GNDA GNDA NE3 W=10u L=5u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM25 net5 net123 GNDA GNDA NE3 W=10u L=5u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM6 VDDA VDDA VDDA VDDA PE3 W=10u L=2u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM5 VDDA VDDA VDDA VDDA PE3 W=10u L=10u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM28 net102 net102 VDDA VDDA PE3 W=10u L=2u M=2.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM0 net7 net7 net102 VDDA PE3 W=10u L=2u M=2.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM23 net6 net6 VDDA VDDA PE3 W=10u L=10u M=8.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM22 net4 net6 VDDA VDDA PE3 W=10u L=10u M=8.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM14 net8 net4 VDDA VDDA PE3 W=10u L=2u M=12.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM4 net1 net4 VDDA VDDA PE3 W=10u L=2u M=10.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM21 RES_BIAS net7 net8 VDDA PE3 W=10u L=1u M=12.0 AD=2.7e-12 AS=3.05e-12 
+ PD=1.054e-05 PS=1.22767e-05 NRD=0.027 NRS=0.027
MM3 OUT2 net7 net1 VDDA PE3 W=10u L=1u M=10.0 AD=2.7e-12 AS=3.12e-12 
+ PD=1.054e-05 PS=1.2624e-05 NRD=0.027 NRS=0.027
MM2 net2 net4 VDDA VDDA PE3 W=10u L=2u M=10.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM1 OUT1 net7 net2 VDDA PE3 W=10u L=1u M=10.0 AD=2.7e-12 AS=3.12e-12 
+ PD=1.054e-05 PS=1.2624e-05 NRD=0.027 NRS=0.027
CC1 net4 net3 $[CMM5T] area=9e-10 perimeter=120.00000u M=8
RR0 net3 RES_BIAS 124.999K $SUB=GNDA $[RPP1K1_3] $W=4u $L=514.1u M=1
XC2 OUT2 GNDA GNDA / mosvc3 W=30u L=30u M=3.0 par1=3.0
XC0 OUT1 GNDA GNDA / mosvc3 W=30u L=30u M=3.0 par1=3.0
.ENDS

************************************************************************
* Library Name: ASKA_BANDGAP
* Cell Name:    bandgap_su
* View Name:    schematic
************************************************************************

.SUBCKT bandgap_su BIAS GNDA OUT VDD3A
*.PININFO BIAS:B GNDA:B OUT:B VDD3A:B
MM29 GNDA GNDA GNDA GNDA NE3 W=10u L=5u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM25 net21 net21 GNDA GNDA NE3 W=1u L=2u M=1.0 AD=4.8e-13 AS=4.8e-13 
+ PD=2.96e-06 PS=2.96e-06 NRD=0.27 NRS=0.27
MM24 VDD3A VDD3A net22 GNDA NE3 W=1u L=2u M=1.0 AD=4.8e-13 AS=4.8e-13 
+ PD=2.96e-06 PS=2.96e-06 NRD=0.27 NRS=0.27
MM23 net22 net22 net21 GNDA NE3 W=1u L=2u M=1.0 AD=4.8e-13 AS=4.8e-13 
+ PD=2.96e-06 PS=2.96e-06 NRD=0.27 NRS=0.27
MM26 GNDA GNDA GNDA GNDA NE3 W=10u L=1u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM17 net12 net21 net7 GNDA NE3 W=10u L=1u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM16 net10 OUT net7 GNDA NE3 W=10u L=1u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM15 net7 net6 GNDA GNDA NE3 W=10u L=1u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM14 net1 net6 GNDA GNDA NE3 W=10u L=1u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM13 OUT net17 GNDA GNDA NE3 W=10u L=1u M=4.0 AD=2.7e-12 AS=3.75e-12 
+ PD=1.054e-05 PS=1.575e-05 NRD=0.027 NRS=0.027
MM11 net3 BIAS net2 GNDA NE3 W=10u L=1u M=4.0 AD=2.7e-12 AS=3.75e-12 
+ PD=1.054e-05 PS=1.575e-05 NRD=0.027 NRS=0.027
MM9 BIAS BIAS net6 GNDA NE3 W=10u L=1u M=4.0 AD=2.7e-12 AS=3.75e-12 
+ PD=1.054e-05 PS=1.575e-05 NRD=0.027 NRS=0.027
MM8 net2 net6 GNDA GNDA NE3 W=10u L=1u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM7 net6 net6 GNDA GNDA NE3 W=10u L=1u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM4 net15 net15 GNDA GNDA NE3 W=10u L=5u M=8.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM2 net17 net15 GNDA GNDA NE3 W=10u L=5u M=8.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM28 A A A VDD3A PE3 W=10u L=5u M=4.0 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 
+ PS=2.096e-05 NRD=0.027 NRS=0.027
MM27 VDD3A VDD3A VDD3A VDD3A PE3 W=10u L=1u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM22 net11 net20 VDD3A VDD3A PE3 W=10u L=5u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM21 net1 net12 net20 VDD3A PE3 W=10u L=5u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM20 net20 net20 VDD3A VDD3A PE3 W=10u L=5u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM19 net12 net10 VDD3A VDD3A PE3 W=10u L=5u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM18 net10 net10 VDD3A VDD3A PE3 W=10u L=5u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM12 OUT net16 VDD3A VDD3A PE3 W=10u L=1u M=16.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM6 net3 net3 net16 VDD3A PE3 W=10u L=1u M=4.0 AD=2.7e-12 AS=3.75e-12 
+ PD=1.054e-05 PS=1.575e-05 NRD=0.027 NRS=0.027
MM1 A net3 net14 VDD3A PE3 W=10u L=1u M=4.0 AD=2.7e-12 AS=3.75e-12 
+ PD=1.054e-05 PS=1.575e-05 NRD=0.027 NRS=0.027
MM0 net16 net16 VDD3A VDD3A PE3 W=10u L=1u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM10 net14 net16 VDD3A VDD3A PE3 W=10u L=1u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM5 net17 net11 A VDD3A PE3 W=10u L=5u M=8.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM3 net15 net23 A VDD3A PE3 W=10u L=5u M=8.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
QQ6 GNDA GNDA net11 QPVC3 1e-10 M=1
QQ5 GNDA GNDA net9 QPVC3 1e-10 M=31
RR11 net5 OUT 200.032K $SUB=GNDA $[RPP1K1_3] $W=4u $L=822.83u M=1
RR10 net8 OUT 200.032K $SUB=GNDA $[RPP1K1_3] $W=4u $L=822.83u M=1
RR8 net23 net5 200.032K $SUB=GNDA $[RPP1K1_3] $W=4u $L=822.83u M=1
RR7 net9 net23 63000 $SUB=GNDA $[RPP1K1_3] $W=8u $L=521.5u M=1
RR6 net11 net8 200.032K $SUB=GNDA $[RPP1K1_3] $W=4u $L=822.83u M=1
CC1 net17 OUT $[CMM5T] area=9e-10 perimeter=120.00000u M=1
.ENDS

************************************************************************
* Library Name: ASKA_BIAS
* Cell Name:    bias
* View Name:    schematic
************************************************************************

.SUBCKT bias BGAP_REF BIAS1 BIAS2 BIAS3 GNDA RES_BIAS VDDA
*.PININFO BGAP_REF:B BIAS1:B BIAS2:B BIAS3:B GNDA:B RES_BIAS:B VDDA:B
XI1 GNDA net2 net1 BIAS3 VDDA / constant_gm
XI2 net2 GNDA BIAS1 BIAS2 RES_BIAS VDDA BGAP_REF / ref_bias
XC0 VDDA GNDA GNDA / mosvc3 W=25.0u L=30u M=26.0 par1=26.0
XI0 net1 GNDA BGAP_REF VDDA / bandgap_su
.ENDS


.SUBCKT mosvc3 G NW SB 
*.PININFO  G:B NW:B SB:B
.ENDS

.SUBCKT ne3i_6 D G S B NW SB 
*.PININFO  D:B G:B S:B B:B NW:B SB:B
.ENDS
