* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : pulse_generator                              *
* Netlisted  : Mon Aug 26 08:47:03 2024                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 LDDN(nedia) nedia2_d dnwtrm(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 1 MN(ne3) nem ndiff(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 2 MP(pe3) pem pdiff(D) p1trm(G) pdiff(S) nwtrm(B)
*.DEVTMPLT 3 NE3I_6() nemi_6 ndiff(D) p1trm(G) ndiff(S) pwitrm(B) dnwtrm(NW) bulk(SB)
*.DEVTMPLT 4 MOSVC3() mosvcm p1trm(G) nwtrm(NW) bulk(SB)
*.DEVTMPLT 5 R(s_res) s_res bulk(POS) bulk(NEG)
*.DEVTMPLT 6 D(p_dnw) p_dnw bulk(POS) nwtrm(NEG)
*.DEVTMPLT 7 D(p_ddnw) p_ddnw bulk(POS) dnwtrm(NEG)
*.DEVTMPLT 8 D(p_dipdnwmv) p_dipwmv pwitrm(POS) dnwtrm(NEG)
*.DEVTMPLT 9 D(p_dnw3) p_dnwm bulk(POS) nwtrm(NEG)
*.DEVTMPLT 10 R(rpp1k1_3) rpp1k1_s p1trm(POS) p1trm(NEG) bulk(SUB)
*.DEVTMPLT 11 R(rpp1k1_3) rpp1k1_n p1trm(POS) p1trm(NEG) nwtrm(SUB)
*.DEVTMPLT 12 C(cmm5t) cmim capm(POS) m4trm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_724654816050                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_724654816050 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_724654816050

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_724654816051                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_724654816051 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_724654816051

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_724654816052                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_724654816052 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_724654816052

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_724654816053                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_724654816053 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_724654816053

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724654816055                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724654816055 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724654816055

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724654816056                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724654816056 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724654816056

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724654816057                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724654816057 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724654816057

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_724654816058                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_724654816058 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_724654816058

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_724654816059                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_724654816059 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_724654816059

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246548160510                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246548160510 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246548160510

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160511                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160511 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246548160511

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160512                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160512 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246548160512

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160513                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160513 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246548160513

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160514                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160514 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246548160514

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160515                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160515 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246548160515

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ND_C_CDNS_7246548160516                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ND_C_CDNS_7246548160516 1 2
** N=2 EP=2 FDC=0
.ends ND_C_CDNS_7246548160516

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246548160517                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246548160517 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246548160517

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160518                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160518 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246548160518

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160519                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160519 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246548160519

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160521                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160521 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246548160521

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246548160522                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246548160522 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246548160522

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160523                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160523 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246548160523

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160524                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160524 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246548160524

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246548160525                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246548160525 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246548160525

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246548160527                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246548160527 1 2
** N=2 EP=2 FDC=0
.ends VIA2_C_CDNS_7246548160527

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160528                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160528 1 2
** N=2 EP=2 FDC=0
.ends VIA1_C_CDNS_7246548160528

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246548160535                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246548160535 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246548160535

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160536                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160536 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246548160536

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_7246548160537                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_7246548160537 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_7246548160537

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160539                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160539 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246548160539

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246548160541                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246548160541 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246548160541

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246548160543                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246548160543 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246548160543

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246548160545                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246548160545 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246548160545

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246548160549                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246548160549 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246548160549

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246548160557                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246548160557 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246548160557

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724654816050                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724654816050 1 2 3
** N=3 EP=3 FDC=4
M0 3 2 1 1 ne3 L=5e-07 W=5e-06 AD=1.35e-12 AS=2.4e-12 PD=5.54e-06 PS=1.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 1 ne3 L=5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=1040 $Y=0 $dt=1
M2 3 2 1 1 ne3 L=5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=2080 $Y=0 $dt=1
M3 1 2 3 1 ne3 L=5e-07 W=5e-06 AD=2.4e-12 AS=1.35e-12 PD=1.096e-05 PS=5.54e-06 $X=3120 $Y=0 $dt=1
.ends ne3_CDNS_724654816050

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nedia_CDNS_724654816051                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nedia_CDNS_724654816051 1 2 3 4
** N=4 EP=4 FDC=1
X0 2 4 3 1 LDDN w=5e-05 l=1.25e-06 adio=1.08602e-09 pdio=0.00013535 extlay=1 $[nedia] $X=-680 $Y=-4850 $dt=0
.ends nedia_CDNS_724654816051

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724654816052                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724654816052 1 2 3
** N=3 EP=3 FDC=4
M0 3 2 1 1 ne3 L=3.5e-07 W=5e-06 AD=1.35e-12 AS=2.4e-12 PD=5.54e-06 PS=1.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 1 ne3 L=3.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=890 $Y=0 $dt=1
M2 3 2 1 1 ne3 L=3.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=1780 $Y=0 $dt=1
M3 1 2 3 1 ne3 L=3.5e-07 W=5e-06 AD=2.4e-12 AS=1.35e-12 PD=1.096e-05 PS=5.54e-06 $X=2670 $Y=0 $dt=1
.ends ne3_CDNS_724654816052

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_724654816053                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_724654816053 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.00010265 W=4e-06 $[rpp1k1_3] $SUB=3 $X=0 $Y=0 $dt=10
.ends rpp1k1_3_CDNS_724654816053

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nedia_CDNS_724654816054                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nedia_CDNS_724654816054 1 2 3 4
** N=4 EP=4 FDC=8
X0 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=-680 $Y=-4850 $dt=0
X1 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=11220 $Y=-4850 $dt=0
X2 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=23120 $Y=-4850 $dt=0
X3 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=35020 $Y=-4850 $dt=0
X4 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=46920 $Y=-4850 $dt=0
X5 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=58820 $Y=-4850 $dt=0
X6 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=70720 $Y=-4850 $dt=0
X7 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=82620 $Y=-4850 $dt=0
.ends nedia_CDNS_724654816054

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724654816055                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724654816055 1 2 3 4
** N=4 EP=4 FDC=2
M0 3 2 1 4 ne3 L=1e-05 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 ne3 L=1e-05 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=10540 $Y=0 $dt=1
.ends ne3_CDNS_724654816055

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724654816056                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724654816056 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=1
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
.ends pe3_CDNS_724654816056

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724654816057                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724654816057 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=2
M0 3 2 1 1 pe3 L=3e-07 W=3e-06 AD=8.1e-13 AS=1.44e-12 PD=3.54e-06 PS=6.96e-06 $X=0 $Y=0 $dt=2
M1 1 2 3 1 pe3 L=3e-07 W=3e-06 AD=1.44e-12 AS=8.1e-13 PD=6.96e-06 PS=3.54e-06 $X=840 $Y=0 $dt=2
.ends pe3_CDNS_724654816057

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_724654816058                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_724654816058 1 2 3
** N=3 EP=3 FDC=1
R0 1 2 L=0.00204354 W=2e-06 $[rpp1k1_3] $SUB=3 $X=-2220 $Y=0 $dt=10
.ends rpp1k1_3_CDNS_724654816058

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160511                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160511 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=1
M0 3 2 1 4 pe3 L=5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
.ends pe3_CDNS_7246548160511

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7246548160512                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7246548160512 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=1e-05 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends ne3_CDNS_7246548160512

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7246548160513                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7246548160513 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=1e-06 W=5e-06 AD=2.4e-12 AS=2.4e-12 PD=1.096e-05 PS=1.096e-05 $X=0 $Y=0 $dt=1
.ends ne3_CDNS_7246548160513

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160514                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160514 1 2 3
*.DEVICECLIMB
** N=3 EP=3 FDC=9
M0 3 2 1 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
M1 1 2 3 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=5540 $Y=0 $dt=2
M2 3 2 1 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=11080 $Y=0 $dt=2
M3 1 2 3 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=16620 $Y=0 $dt=2
M4 3 2 1 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=22160 $Y=0 $dt=2
M5 1 2 3 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=27700 $Y=0 $dt=2
M6 3 2 1 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=33240 $Y=0 $dt=2
M7 1 2 3 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=38780 $Y=0 $dt=2
M8 3 2 1 1 pe3 L=5e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=44320 $Y=0 $dt=2
.ends pe3_CDNS_7246548160514

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7246548160515                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7246548160515 1 2 3
** N=3 EP=3 FDC=1
R0 1 2 L=1e-05 W=2e-06 $[rpp1k1_3] $SUB=3 $X=0 $Y=0 $dt=10
.ends rpp1k1_3_CDNS_7246548160515

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7246548160516                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7246548160516 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
R0 2 1 L=0.00016435 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=11
.ends rpp1k1_3_CDNS_7246548160516

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7246548160517                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7246548160517 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.00041122 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=10
.ends rpp1k1_3_CDNS_7246548160517

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7246548160518                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7246548160518 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=3.5e-07 W=2e-06 AD=9.6e-13 AS=9.6e-13 PD=4.96e-06 PS=4.96e-06 $X=0 $Y=0 $dt=1
.ends ne3_CDNS_7246548160518

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246548160548                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246548160548 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246548160548

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X1 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7246548160548 $T=660 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7246548160548 $T=660 1500 0 0 $X=0 $Y=1000
X2 1 VIATP_C_CDNS_7246548160548 $T=660 2500 0 0 $X=0 $Y=2000
X3 1 VIATP_C_CDNS_7246548160548 $T=660 3500 0 0 $X=0 $Y=3000
X4 1 VIATP_C_CDNS_7246548160548 $T=660 4500 0 0 $X=0 $Y=4000
.ends MASCO__X1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246548160547                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246548160547 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246548160547

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X2 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7246548160547 $T=790 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7246548160547 $T=790 1500 0 0 $X=0 $Y=1000
X2 1 VIATP_C_CDNS_7246548160547 $T=790 2500 0 0 $X=0 $Y=2000
X3 1 VIATP_C_CDNS_7246548160547 $T=790 3500 0 0 $X=0 $Y=3000
X4 1 VIATP_C_CDNS_7246548160547 $T=790 4500 0 0 $X=0 $Y=4000
.ends MASCO__X2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246548160546                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246548160546 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246548160546

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X5                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X5 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7246548160546 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7246548160546 $T=500 1500 0 0 $X=0 $Y=1000
X2 1 VIATP_C_CDNS_7246548160546 $T=500 2500 0 0 $X=0 $Y=2000
X3 1 VIATP_C_CDNS_7246548160546 $T=500 3500 0 0 $X=0 $Y=3000
X4 1 VIATP_C_CDNS_7246548160546 $T=500 4500 0 0 $X=0 $Y=4000
.ends MASCO__X5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y6                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y6 1
** N=1 EP=1 FDC=0
X0 1 MASCO__X5 $T=0 0 0 0 $X=0 $Y=0
X1 1 MASCO__X5 $T=2000 0 0 0 $X=2000 $Y=0
X2 1 MASCO__X5 $T=4000 0 0 0 $X=4000 $Y=0
X3 1 MASCO__X5 $T=6000 0 0 0 $X=6000 $Y=0
X4 1 MASCO__X5 $T=8000 0 0 0 $X=8000 $Y=0
X5 1 MASCO__X5 $T=10000 0 0 0 $X=10000 $Y=0
X6 1 MASCO__X5 $T=12000 0 0 0 $X=12000 $Y=0
X7 1 MASCO__X5 $T=14000 0 0 0 $X=14000 $Y=0
X8 1 MASCO__X5 $T=16000 0 0 0 $X=16000 $Y=0
.ends MASCO__Y6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X4                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X4 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7246548160546 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7246548160546 $T=500 2500 0 0 $X=0 $Y=2000
X2 1 VIATP_C_CDNS_7246548160546 $T=500 4500 0 0 $X=0 $Y=4000
X3 1 VIATP_C_CDNS_7246548160546 $T=500 6500 0 0 $X=0 $Y=6000
X4 1 VIATP_C_CDNS_7246548160546 $T=500 8500 0 0 $X=0 $Y=8000
X5 1 VIATP_C_CDNS_7246548160546 $T=500 10500 0 0 $X=0 $Y=10000
X6 1 VIATP_C_CDNS_7246548160546 $T=500 12500 0 0 $X=0 $Y=12000
X7 1 VIATP_C_CDNS_7246548160546 $T=500 14500 0 0 $X=0 $Y=14000
X8 1 VIATP_C_CDNS_7246548160546 $T=500 16500 0 0 $X=0 $Y=16000
X9 1 VIATP_C_CDNS_7246548160546 $T=500 18500 0 0 $X=0 $Y=18000
X10 1 VIATP_C_CDNS_7246548160546 $T=500 20500 0 0 $X=0 $Y=20000
X11 1 VIATP_C_CDNS_7246548160546 $T=500 22500 0 0 $X=0 $Y=22000
.ends MASCO__X4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y7                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y7 1
** N=1 EP=1 FDC=0
X0 1 MASCO__X4 $T=0 0 0 0 $X=0 $Y=0
X1 1 MASCO__X4 $T=2000 0 0 0 $X=2000 $Y=0
X2 1 MASCO__X4 $T=4000 0 0 0 $X=4000 $Y=0
X3 1 MASCO__X4 $T=6000 0 0 0 $X=6000 $Y=0
X4 1 MASCO__X4 $T=8000 0 0 0 $X=8000 $Y=0
X5 1 MASCO__X4 $T=10000 0 0 0 $X=10000 $Y=0
X6 1 MASCO__X4 $T=12000 0 0 0 $X=12000 $Y=0
.ends MASCO__Y7

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X3                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X3 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7246548160546 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7246548160546 $T=500 2500 0 0 $X=0 $Y=2000
X2 1 VIATP_C_CDNS_7246548160546 $T=500 4500 0 0 $X=0 $Y=4000
X3 1 VIATP_C_CDNS_7246548160546 $T=500 6500 0 0 $X=0 $Y=6000
X4 1 VIATP_C_CDNS_7246548160546 $T=500 8500 0 0 $X=0 $Y=8000
X5 1 VIATP_C_CDNS_7246548160546 $T=500 10500 0 0 $X=0 $Y=10000
X6 1 VIATP_C_CDNS_7246548160546 $T=500 12500 0 0 $X=0 $Y=12000
X7 1 VIATP_C_CDNS_7246548160546 $T=500 14500 0 0 $X=0 $Y=14000
X8 1 VIATP_C_CDNS_7246548160546 $T=500 16500 0 0 $X=0 $Y=16000
X9 1 VIATP_C_CDNS_7246548160546 $T=500 18500 0 0 $X=0 $Y=18000
X10 1 VIATP_C_CDNS_7246548160546 $T=500 20500 0 0 $X=0 $Y=20000
.ends MASCO__X3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y8                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y8 1
** N=1 EP=1 FDC=0
X0 1 MASCO__X3 $T=0 0 0 0 $X=0 $Y=0
X1 1 MASCO__X3 $T=2000 0 0 0 $X=2000 $Y=0
X2 1 MASCO__X3 $T=4000 0 0 0 $X=4000 $Y=0
X3 1 MASCO__X3 $T=6000 0 0 0 $X=6000 $Y=0
X4 1 MASCO__X3 $T=8000 0 0 0 $X=8000 $Y=0
X5 1 MASCO__X3 $T=10000 0 0 0 $X=10000 $Y=0
X6 1 MASCO__X3 $T=12000 0 0 0 $X=12000 $Y=0
.ends MASCO__Y8

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246548160544                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246548160544 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246548160544

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y9                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y9 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7246548160544 $T=500 530 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7246548160544 $T=1500 530 0 0 $X=1000 $Y=0
X2 1 VIATP_C_CDNS_7246548160544 $T=2500 530 0 0 $X=2000 $Y=0
X3 1 VIATP_C_CDNS_7246548160544 $T=3500 530 0 0 $X=3000 $Y=0
X4 1 VIATP_C_CDNS_7246548160544 $T=4500 530 0 0 $X=4000 $Y=0
X5 1 VIATP_C_CDNS_7246548160544 $T=5500 530 0 0 $X=5000 $Y=0
X6 1 VIATP_C_CDNS_7246548160544 $T=6500 530 0 0 $X=6000 $Y=0
X7 1 VIATP_C_CDNS_7246548160544 $T=7500 530 0 0 $X=7000 $Y=0
X8 1 VIATP_C_CDNS_7246548160544 $T=8500 530 0 0 $X=8000 $Y=0
X9 1 VIATP_C_CDNS_7246548160544 $T=9500 530 0 0 $X=9000 $Y=0
X10 1 VIATP_C_CDNS_7246548160544 $T=10500 530 0 0 $X=10000 $Y=0
.ends MASCO__Y9

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: current_source_gm_10_en_r                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt current_source_gm_10_en_r 1 2 3 4 5 6 7 8 9 10
+ 11
*.DEVICECLIMB
** N=27 EP=11 FDC=197
X0 6 VIA3_C_CDNS_724654816050 $T=98240 32160 0 0 $X=97490 $Y=31410
X1 12 VIA1_C_CDNS_724654816055 $T=7790 61030 0 0 $X=7390 $Y=60320
X2 4 VIA1_C_CDNS_724654816055 $T=18330 62810 0 0 $X=17930 $Y=62100
X3 12 VIA1_C_CDNS_724654816055 $T=28870 61030 0 0 $X=28470 $Y=60320
X4 13 VIA1_C_CDNS_724654816055 $T=33575 62810 0 0 $X=33175 $Y=62100
X5 14 VIA1_C_CDNS_724654816055 $T=44115 61030 0 0 $X=43715 $Y=60320
X6 13 VIA1_C_CDNS_724654816055 $T=54655 62810 0 0 $X=54255 $Y=62100
X7 15 VIA1_C_CDNS_724654816055 $T=59300 62950 0 0 $X=58900 $Y=62240
X8 16 VIA1_C_CDNS_724654816055 $T=69840 61110 0 0 $X=69440 $Y=60400
X9 15 VIA1_C_CDNS_724654816055 $T=80380 62950 0 0 $X=79980 $Y=62240
X10 17 VIA1_C_CDNS_724654816055 $T=106545 17830 0 0 $X=106145 $Y=17120
X11 18 VIA1_C_CDNS_724654816055 $T=106545 45950 0 0 $X=106145 $Y=45240
X12 17 VIA1_C_CDNS_724654816055 $T=117625 17830 0 0 $X=117225 $Y=17120
X13 18 VIA1_C_CDNS_724654816055 $T=117625 45950 0 0 $X=117225 $Y=45240
X14 17 VIA1_C_CDNS_724654816055 $T=128705 17830 0 0 $X=128305 $Y=17120
X15 18 VIA1_C_CDNS_724654816055 $T=128705 45950 0 0 $X=128305 $Y=45240
X16 17 VIA1_C_CDNS_724654816055 $T=139785 17830 0 0 $X=139385 $Y=17120
X17 18 VIA1_C_CDNS_724654816055 $T=139785 45950 0 0 $X=139385 $Y=45240
X18 17 VIA1_C_CDNS_724654816055 $T=150865 17830 0 0 $X=150465 $Y=17120
X19 18 VIA1_C_CDNS_724654816055 $T=150865 45950 0 0 $X=150465 $Y=45240
X20 18 VIA1_C_CDNS_724654816055 $T=160825 16050 0 0 $X=160425 $Y=15340
X21 17 VIA1_C_CDNS_724654816055 $T=160825 47730 0 0 $X=160425 $Y=47020
X22 18 VIA1_C_CDNS_724654816055 $T=171905 16050 0 0 $X=171505 $Y=15340
X23 17 VIA1_C_CDNS_724654816055 $T=171905 47730 0 0 $X=171505 $Y=47020
X24 18 VIA1_C_CDNS_724654816055 $T=182985 16050 0 0 $X=182585 $Y=15340
X25 17 VIA1_C_CDNS_724654816055 $T=182985 47730 0 0 $X=182585 $Y=47020
X26 18 VIA1_C_CDNS_724654816055 $T=194065 16050 0 0 $X=193665 $Y=15340
X27 17 VIA1_C_CDNS_724654816055 $T=194065 47730 0 0 $X=193665 $Y=47020
X28 18 VIA1_C_CDNS_724654816055 $T=205145 16050 0 0 $X=204745 $Y=15340
X29 17 VIA1_C_CDNS_724654816055 $T=205145 47730 0 0 $X=204745 $Y=47020
X30 1 VIA1_C_CDNS_724654816056 $T=247850 19860 0 0 $X=247710 $Y=18890
X31 19 VIA1_C_CDNS_724654816056 $T=248890 17580 0 0 $X=248750 $Y=16610
X32 1 VIA1_C_CDNS_724654816056 $T=249930 19860 0 0 $X=249790 $Y=18890
X33 19 VIA1_C_CDNS_724654816056 $T=250970 17580 0 0 $X=250830 $Y=16610
X34 1 VIA1_C_CDNS_724654816056 $T=252010 19860 0 0 $X=251870 $Y=18890
X35 12 VIA1_C_CDNS_724654816057 $T=33660 31900 0 0 $X=33260 $Y=31710
X36 12 VIA1_C_CDNS_724654816057 $T=44900 31900 0 0 $X=44500 $Y=31710
X37 12 VIA1_C_CDNS_724654816057 $T=56140 31900 0 0 $X=55740 $Y=31710
X38 14 VIA1_C_CDNS_724654816057 $T=63465 83370 0 0 $X=63065 $Y=83180
X39 14 VIA1_C_CDNS_724654816057 $T=65705 83370 0 0 $X=65305 $Y=83180
X40 14 VIA1_C_CDNS_724654816057 $T=67945 83370 0 0 $X=67545 $Y=83180
X41 14 VIA1_C_CDNS_724654816057 $T=70185 83370 0 0 $X=69785 $Y=83180
X42 14 VIA1_C_CDNS_724654816057 $T=72425 83370 0 0 $X=72025 $Y=83180
X43 17 VIA1_C_CDNS_724654816057 $T=117900 81120 0 0 $X=117500 $Y=80930
X44 18 VIA1_C_CDNS_724654816057 $T=119550 81900 0 0 $X=119150 $Y=81710
X45 16 VIA1_C_CDNS_724654816057 $T=122400 137545 0 0 $X=122000 $Y=137355
X46 17 VIA1_C_CDNS_724654816057 $T=124680 81120 0 0 $X=124280 $Y=80930
X47 18 VIA1_C_CDNS_724654816057 $T=125360 81900 0 0 $X=124960 $Y=81710
X48 16 VIA1_C_CDNS_724654816057 $T=128640 137545 0 0 $X=128240 $Y=137355
X49 17 VIA1_C_CDNS_724654816057 $T=130380 81120 0 0 $X=129980 $Y=80930
X50 18 VIA1_C_CDNS_724654816057 $T=132030 81900 0 0 $X=131630 $Y=81710
X51 16 VIA1_C_CDNS_724654816057 $T=134880 137545 0 0 $X=134480 $Y=137355
X52 17 VIA1_C_CDNS_724654816057 $T=137160 81120 0 0 $X=136760 $Y=80930
X53 18 VIA1_C_CDNS_724654816057 $T=137840 81900 0 0 $X=137440 $Y=81710
X54 16 VIA1_C_CDNS_724654816057 $T=141120 137545 0 0 $X=140720 $Y=137355
X55 17 VIA1_C_CDNS_724654816057 $T=142860 81120 0 0 $X=142460 $Y=80930
X56 18 VIA1_C_CDNS_724654816057 $T=144510 81900 0 0 $X=144110 $Y=81710
X57 16 VIA1_C_CDNS_724654816057 $T=147360 137545 0 0 $X=146960 $Y=137355
X58 17 VIA1_C_CDNS_724654816057 $T=149640 81120 0 0 $X=149240 $Y=80930
X59 18 VIA1_C_CDNS_724654816057 $T=150320 81900 0 0 $X=149920 $Y=81710
X60 16 VIA1_C_CDNS_724654816057 $T=153600 137545 0 0 $X=153200 $Y=137355
X61 17 VIA1_C_CDNS_724654816057 $T=155340 81120 0 0 $X=154940 $Y=80930
X62 18 VIA1_C_CDNS_724654816057 $T=156990 81900 0 0 $X=156590 $Y=81710
X63 16 VIA1_C_CDNS_724654816057 $T=159840 137545 0 0 $X=159440 $Y=137355
X64 17 VIA1_C_CDNS_724654816057 $T=162120 81120 0 0 $X=161720 $Y=80930
X65 18 VIA1_C_CDNS_724654816057 $T=162800 81900 0 0 $X=162400 $Y=81710
X66 16 VIA1_C_CDNS_724654816057 $T=166080 137545 0 0 $X=165680 $Y=137355
X67 17 VIA1_C_CDNS_724654816057 $T=167820 81120 0 0 $X=167420 $Y=80930
X68 18 VIA1_C_CDNS_724654816057 $T=169470 81900 0 0 $X=169070 $Y=81710
X69 16 VIA1_C_CDNS_724654816057 $T=172320 137545 0 0 $X=171920 $Y=137355
X70 17 VIA1_C_CDNS_724654816057 $T=174600 81120 0 0 $X=174200 $Y=80930
X71 18 VIA1_C_CDNS_724654816057 $T=175280 81900 0 0 $X=174880 $Y=81710
X72 16 VIA1_C_CDNS_724654816057 $T=178560 137545 0 0 $X=178160 $Y=137355
X73 17 VIA1_C_CDNS_724654816057 $T=180300 81120 0 0 $X=179900 $Y=80930
X74 18 VIA1_C_CDNS_724654816057 $T=181950 81900 0 0 $X=181550 $Y=81710
X75 16 VIA1_C_CDNS_724654816057 $T=184800 137545 0 0 $X=184400 $Y=137355
X76 17 VIA1_C_CDNS_724654816057 $T=187080 81120 0 0 $X=186680 $Y=80930
X77 18 VIA1_C_CDNS_724654816057 $T=187760 81900 0 0 $X=187360 $Y=81710
X78 16 VIA1_C_CDNS_724654816057 $T=191040 137545 0 0 $X=190640 $Y=137355
X79 17 VIA1_C_CDNS_724654816057 $T=192780 81120 0 0 $X=192380 $Y=80930
X80 18 VIA1_C_CDNS_724654816057 $T=194430 81900 0 0 $X=194030 $Y=81710
X81 16 VIA1_C_CDNS_724654816057 $T=197280 137545 0 0 $X=196880 $Y=137355
X82 17 VIA1_C_CDNS_724654816057 $T=199560 81120 0 0 $X=199160 $Y=80930
X83 18 VIA1_C_CDNS_724654816057 $T=200240 81900 0 0 $X=199840 $Y=81710
X84 20 VIA1_C_CDNS_724654816057 $T=248180 27500 0 0 $X=247780 $Y=27310
X85 20 VIA1_C_CDNS_724654816057 $T=249410 27500 0 0 $X=249010 $Y=27310
X86 20 VIA1_C_CDNS_724654816057 $T=250450 27500 0 0 $X=250050 $Y=27310
X87 20 VIA1_C_CDNS_724654816057 $T=251680 27500 0 0 $X=251280 $Y=27310
X88 12 VIA2_C_CDNS_724654816058 $T=8380 17610 0 0 $X=7410 $Y=16950
X89 12 VIA2_C_CDNS_724654816058 $T=8380 49670 0 0 $X=7410 $Y=49010
X90 13 VIA2_C_CDNS_724654816058 $T=10660 15770 0 0 $X=9690 $Y=15110
X91 13 VIA2_C_CDNS_724654816058 $T=10660 47830 0 0 $X=9690 $Y=47170
X92 15 VIA2_C_CDNS_724654816058 $T=12940 13930 0 0 $X=11970 $Y=13270
X93 15 VIA2_C_CDNS_724654816058 $T=12940 45990 0 0 $X=11970 $Y=45330
X94 13 VIA2_C_CDNS_724654816058 $T=76860 15770 0 0 $X=75890 $Y=15110
X95 13 VIA2_C_CDNS_724654816058 $T=76860 47830 0 0 $X=75890 $Y=47170
X96 15 VIA2_C_CDNS_724654816058 $T=79200 13930 0 0 $X=78230 $Y=13270
X97 15 VIA2_C_CDNS_724654816058 $T=79200 45990 0 0 $X=78230 $Y=45330
X98 12 VIA2_C_CDNS_724654816058 $T=81540 17610 0 0 $X=80570 $Y=16950
X99 12 VIA2_C_CDNS_724654816058 $T=81540 49670 0 0 $X=80570 $Y=49010
X100 20 VIA2_C_CDNS_724654816058 $T=102350 65860 0 0 $X=101380 $Y=65200
X101 20 VIA2_C_CDNS_724654816058 $T=102350 98940 0 0 $X=101380 $Y=98280
X102 16 VIA2_C_CDNS_724654816058 $T=104030 116805 0 0 $X=103060 $Y=116145
X103 16 VIA2_C_CDNS_724654816058 $T=104030 158145 0 0 $X=103060 $Y=157485
X104 21 VIA2_C_CDNS_724654816058 $T=104630 64080 0 0 $X=103660 $Y=63420
X105 21 VIA2_C_CDNS_724654816058 $T=104630 97160 0 0 $X=103660 $Y=96500
X106 17 VIA2_C_CDNS_724654816058 $T=106310 120365 0 0 $X=105340 $Y=119705
X107 17 VIA2_C_CDNS_724654816058 $T=106310 152805 0 0 $X=105340 $Y=152145
X108 22 VIA2_C_CDNS_724654816058 $T=106910 67640 0 0 $X=105940 $Y=66980
X109 22 VIA2_C_CDNS_724654816058 $T=106910 95380 0 0 $X=105940 $Y=94720
X110 22 VIA2_C_CDNS_724654816058 $T=108590 118585 0 0 $X=107620 $Y=117925
X111 22 VIA2_C_CDNS_724654816058 $T=108590 156365 0 0 $X=107620 $Y=155705
X112 2 VIA2_C_CDNS_724654816058 $T=110870 123925 0 0 $X=109900 $Y=123265
X113 2 VIA2_C_CDNS_724654816058 $T=110870 151025 0 0 $X=109900 $Y=150365
X114 2 VIA2_C_CDNS_724654816058 $T=208810 123925 0 0 $X=207840 $Y=123265
X115 2 VIA2_C_CDNS_724654816058 $T=208810 151025 0 0 $X=207840 $Y=150365
X116 22 VIA2_C_CDNS_724654816058 $T=211090 67640 0 0 $X=210120 $Y=66980
X117 22 VIA2_C_CDNS_724654816058 $T=211090 95380 0 0 $X=210120 $Y=94720
X118 22 VIA2_C_CDNS_724654816058 $T=211090 118585 0 0 $X=210120 $Y=117925
X119 22 VIA2_C_CDNS_724654816058 $T=211090 156365 0 0 $X=210120 $Y=155705
X120 20 VIA2_C_CDNS_724654816058 $T=213370 65860 0 0 $X=212400 $Y=65200
X121 20 VIA2_C_CDNS_724654816058 $T=213370 98940 0 0 $X=212400 $Y=98280
X122 18 VIA2_C_CDNS_724654816058 $T=213370 122145 0 0 $X=212400 $Y=121485
X123 18 VIA2_C_CDNS_724654816058 $T=213370 154585 0 0 $X=212400 $Y=153925
X124 21 VIA2_C_CDNS_724654816058 $T=215650 64080 0 0 $X=214680 $Y=63420
X125 21 VIA2_C_CDNS_724654816058 $T=215650 97160 0 0 $X=214680 $Y=96500
X126 16 VIA2_C_CDNS_724654816058 $T=215650 116805 0 0 $X=214680 $Y=116145
X127 16 VIA2_C_CDNS_724654816058 $T=215650 158145 0 0 $X=214680 $Y=157485
X128 20 VIA2_C_CDNS_724654816058 $T=227815 16050 0 0 $X=226845 $Y=15390
X129 20 VIA2_C_CDNS_724654816058 $T=227815 37420 0 0 $X=226845 $Y=36760
X130 21 VIA2_C_CDNS_724654816058 $T=239775 17830 0 0 $X=238805 $Y=17170
X131 21 VIA2_C_CDNS_724654816058 $T=239775 35640 0 0 $X=238805 $Y=34980
X132 13 VIA2_C_CDNS_724654816059 $T=44040 62810 0 0 $X=41990 $Y=62060
X133 15 VIA2_C_CDNS_724654816059 $T=78860 62950 0 0 $X=76810 $Y=62200
X134 23 VIA2_C_CDNS_724654816059 $T=311195 26360 0 0 $X=309145 $Y=25610
X135 9 VIA2_C_CDNS_724654816059 $T=315635 26360 0 0 $X=313585 $Y=25610
X136 23 VIA2_C_CDNS_724654816059 $T=324920 82035 0 0 $X=322870 $Y=81285
X137 12 VIA2_C_CDNS_7246548160510 $T=8380 31900 0 0 $X=7410 $Y=31760
X138 12 VIA2_C_CDNS_7246548160510 $T=81540 31900 0 0 $X=80570 $Y=31760
X139 16 VIA2_C_CDNS_7246548160510 $T=104030 137545 0 0 $X=103060 $Y=137405
X140 16 VIA2_C_CDNS_7246548160510 $T=215650 137545 0 0 $X=214680 $Y=137405
X141 1 VIA1_C_CDNS_7246548160511 $T=15280 19450 0 0 $X=14310 $Y=18790
X142 1 VIA1_C_CDNS_7246548160511 $T=15280 44150 0 0 $X=14310 $Y=43490
X143 1 VIA1_C_CDNS_7246548160511 $T=74520 19450 0 0 $X=73550 $Y=18790
X144 1 VIA1_C_CDNS_7246548160511 $T=74520 44150 0 0 $X=73550 $Y=43490
X145 1 VIA1_C_CDNS_7246548160511 $T=230095 19610 0 0 $X=229125 $Y=18950
X146 1 VIA1_C_CDNS_7246548160511 $T=230095 33860 0 0 $X=229125 $Y=33200
X147 1 VIA1_C_CDNS_7246548160511 $T=237495 19610 0 0 $X=236525 $Y=18950
X148 1 VIA1_C_CDNS_7246548160511 $T=237495 33860 0 0 $X=236525 $Y=33200
X149 21 VIA1_C_CDNS_7246548160512 $T=201995 64080 0 0 $X=201545 $Y=63680
X150 20 VIA1_C_CDNS_7246548160512 $T=201995 98940 0 0 $X=201545 $Y=98540
X151 22 VIA1_C_CDNS_7246548160513 $T=115670 67640 0 0 $X=115480 $Y=66980
X152 22 VIA1_C_CDNS_7246548160513 $T=115670 95380 0 0 $X=115480 $Y=94720
X153 20 VIA1_C_CDNS_7246548160513 $T=121210 65860 0 0 $X=121020 $Y=65200
X154 21 VIA1_C_CDNS_7246548160513 $T=121210 97160 0 0 $X=121020 $Y=96500
X155 22 VIA1_C_CDNS_7246548160513 $T=121910 67640 0 0 $X=121720 $Y=66980
X156 22 VIA1_C_CDNS_7246548160513 $T=121910 95380 0 0 $X=121720 $Y=94720
X157 21 VIA1_C_CDNS_7246548160513 $T=127450 64080 0 0 $X=127260 $Y=63420
X158 20 VIA1_C_CDNS_7246548160513 $T=127450 98940 0 0 $X=127260 $Y=98280
X159 22 VIA1_C_CDNS_7246548160513 $T=128150 67640 0 0 $X=127960 $Y=66980
X160 22 VIA1_C_CDNS_7246548160513 $T=128150 95380 0 0 $X=127960 $Y=94720
X161 20 VIA1_C_CDNS_7246548160513 $T=133690 65860 0 0 $X=133500 $Y=65200
X162 21 VIA1_C_CDNS_7246548160513 $T=133690 97160 0 0 $X=133500 $Y=96500
X163 22 VIA1_C_CDNS_7246548160513 $T=134390 67640 0 0 $X=134200 $Y=66980
X164 22 VIA1_C_CDNS_7246548160513 $T=134390 95380 0 0 $X=134200 $Y=94720
X165 21 VIA1_C_CDNS_7246548160513 $T=139930 64080 0 0 $X=139740 $Y=63420
X166 20 VIA1_C_CDNS_7246548160513 $T=139930 98940 0 0 $X=139740 $Y=98280
X167 22 VIA1_C_CDNS_7246548160513 $T=140630 67640 0 0 $X=140440 $Y=66980
X168 22 VIA1_C_CDNS_7246548160513 $T=140630 95380 0 0 $X=140440 $Y=94720
X169 20 VIA1_C_CDNS_7246548160513 $T=146170 65860 0 0 $X=145980 $Y=65200
X170 21 VIA1_C_CDNS_7246548160513 $T=146170 97160 0 0 $X=145980 $Y=96500
X171 22 VIA1_C_CDNS_7246548160513 $T=146870 67640 0 0 $X=146680 $Y=66980
X172 22 VIA1_C_CDNS_7246548160513 $T=146870 95380 0 0 $X=146680 $Y=94720
X173 21 VIA1_C_CDNS_7246548160513 $T=152410 64080 0 0 $X=152220 $Y=63420
X174 20 VIA1_C_CDNS_7246548160513 $T=152410 98940 0 0 $X=152220 $Y=98280
X175 22 VIA1_C_CDNS_7246548160513 $T=153110 67640 0 0 $X=152920 $Y=66980
X176 22 VIA1_C_CDNS_7246548160513 $T=153110 95380 0 0 $X=152920 $Y=94720
X177 20 VIA1_C_CDNS_7246548160513 $T=158650 65860 0 0 $X=158460 $Y=65200
X178 21 VIA1_C_CDNS_7246548160513 $T=158650 97160 0 0 $X=158460 $Y=96500
X179 22 VIA1_C_CDNS_7246548160513 $T=159350 67640 0 0 $X=159160 $Y=66980
X180 22 VIA1_C_CDNS_7246548160513 $T=159350 95380 0 0 $X=159160 $Y=94720
X181 21 VIA1_C_CDNS_7246548160513 $T=164890 64080 0 0 $X=164700 $Y=63420
X182 20 VIA1_C_CDNS_7246548160513 $T=164890 98940 0 0 $X=164700 $Y=98280
X183 22 VIA1_C_CDNS_7246548160513 $T=165590 67640 0 0 $X=165400 $Y=66980
X184 22 VIA1_C_CDNS_7246548160513 $T=165590 95380 0 0 $X=165400 $Y=94720
X185 20 VIA1_C_CDNS_7246548160513 $T=171130 65860 0 0 $X=170940 $Y=65200
X186 21 VIA1_C_CDNS_7246548160513 $T=171130 97160 0 0 $X=170940 $Y=96500
X187 22 VIA1_C_CDNS_7246548160513 $T=171830 67640 0 0 $X=171640 $Y=66980
X188 22 VIA1_C_CDNS_7246548160513 $T=171830 95380 0 0 $X=171640 $Y=94720
X189 21 VIA1_C_CDNS_7246548160513 $T=177370 64080 0 0 $X=177180 $Y=63420
X190 20 VIA1_C_CDNS_7246548160513 $T=177370 98940 0 0 $X=177180 $Y=98280
X191 22 VIA1_C_CDNS_7246548160513 $T=178070 67640 0 0 $X=177880 $Y=66980
X192 22 VIA1_C_CDNS_7246548160513 $T=178070 95380 0 0 $X=177880 $Y=94720
X193 20 VIA1_C_CDNS_7246548160513 $T=183610 65860 0 0 $X=183420 $Y=65200
X194 21 VIA1_C_CDNS_7246548160513 $T=183610 97160 0 0 $X=183420 $Y=96500
X195 22 VIA1_C_CDNS_7246548160513 $T=184310 67640 0 0 $X=184120 $Y=66980
X196 22 VIA1_C_CDNS_7246548160513 $T=184310 95380 0 0 $X=184120 $Y=94720
X197 21 VIA1_C_CDNS_7246548160513 $T=189850 64080 0 0 $X=189660 $Y=63420
X198 20 VIA1_C_CDNS_7246548160513 $T=189850 98940 0 0 $X=189660 $Y=98280
X199 22 VIA1_C_CDNS_7246548160513 $T=190550 67640 0 0 $X=190360 $Y=66980
X200 22 VIA1_C_CDNS_7246548160513 $T=190550 95380 0 0 $X=190360 $Y=94720
X201 20 VIA1_C_CDNS_7246548160513 $T=196090 65860 0 0 $X=195900 $Y=65200
X202 21 VIA1_C_CDNS_7246548160513 $T=196090 97160 0 0 $X=195900 $Y=96500
X203 22 VIA1_C_CDNS_7246548160513 $T=196790 67640 0 0 $X=196600 $Y=66980
X204 22 VIA1_C_CDNS_7246548160513 $T=196790 95380 0 0 $X=196600 $Y=94720
X205 1 VIA1_C_CDNS_7246548160514 $T=17150 19450 0 0 $X=17010 $Y=18740
X206 1 VIA1_C_CDNS_7246548160514 $T=17150 44150 0 0 $X=17010 $Y=43440
X207 1 VIA1_C_CDNS_7246548160514 $T=27690 19450 0 0 $X=27550 $Y=18740
X208 1 VIA1_C_CDNS_7246548160514 $T=27690 44150 0 0 $X=27550 $Y=43440
X209 1 VIA1_C_CDNS_7246548160514 $T=28390 19450 0 0 $X=28250 $Y=18740
X210 1 VIA1_C_CDNS_7246548160514 $T=28390 44150 0 0 $X=28250 $Y=43440
X211 15 VIA1_C_CDNS_7246548160514 $T=38930 13930 0 0 $X=38790 $Y=13220
X212 15 VIA1_C_CDNS_7246548160514 $T=38930 45990 0 0 $X=38790 $Y=45280
X213 1 VIA1_C_CDNS_7246548160514 $T=39630 19450 0 0 $X=39490 $Y=18740
X214 1 VIA1_C_CDNS_7246548160514 $T=39630 44150 0 0 $X=39490 $Y=43440
X215 12 VIA1_C_CDNS_7246548160514 $T=50170 17610 0 0 $X=50030 $Y=16900
X216 12 VIA1_C_CDNS_7246548160514 $T=50170 49670 0 0 $X=50030 $Y=48960
X217 1 VIA1_C_CDNS_7246548160514 $T=50870 19450 0 0 $X=50730 $Y=18740
X218 1 VIA1_C_CDNS_7246548160514 $T=50870 44150 0 0 $X=50730 $Y=43440
X219 13 VIA1_C_CDNS_7246548160514 $T=61410 15770 0 0 $X=61270 $Y=15060
X220 13 VIA1_C_CDNS_7246548160514 $T=61410 47830 0 0 $X=61270 $Y=47120
X221 1 VIA1_C_CDNS_7246548160514 $T=62110 19450 0 0 $X=61970 $Y=18740
X222 1 VIA1_C_CDNS_7246548160514 $T=62110 44150 0 0 $X=61970 $Y=43440
X223 19 VIA1_C_CDNS_7246548160514 $T=62695 100410 0 0 $X=62555 $Y=99700
X224 2 VIA1_C_CDNS_7246548160514 $T=64235 96850 0 0 $X=64095 $Y=96140
X225 19 VIA1_C_CDNS_7246548160514 $T=64935 100410 0 0 $X=64795 $Y=99700
X226 2 VIA1_C_CDNS_7246548160514 $T=66475 96850 0 0 $X=66335 $Y=96140
X227 14 VIA1_C_CDNS_7246548160514 $T=67175 98630 0 0 $X=67035 $Y=97920
X228 2 VIA1_C_CDNS_7246548160514 $T=68715 96850 0 0 $X=68575 $Y=96140
X229 19 VIA1_C_CDNS_7246548160514 $T=69415 100410 0 0 $X=69275 $Y=99700
X230 2 VIA1_C_CDNS_7246548160514 $T=70955 96850 0 0 $X=70815 $Y=96140
X231 19 VIA1_C_CDNS_7246548160514 $T=71655 100410 0 0 $X=71515 $Y=99700
X232 1 VIA1_C_CDNS_7246548160514 $T=72650 19450 0 0 $X=72510 $Y=18740
X233 1 VIA1_C_CDNS_7246548160514 $T=72650 44150 0 0 $X=72510 $Y=43440
X234 2 VIA1_C_CDNS_7246548160514 $T=73195 96850 0 0 $X=73055 $Y=96140
X235 2 VIA1_C_CDNS_7246548160514 $T=113390 123925 0 0 $X=113250 $Y=123215
X236 2 VIA1_C_CDNS_7246548160514 $T=113390 151025 0 0 $X=113250 $Y=150315
X237 2 VIA1_C_CDNS_7246548160514 $T=118930 123925 0 0 $X=118790 $Y=123215
X238 2 VIA1_C_CDNS_7246548160514 $T=118930 151025 0 0 $X=118790 $Y=150315
X239 2 VIA1_C_CDNS_7246548160514 $T=119630 123925 0 0 $X=119490 $Y=123215
X240 2 VIA1_C_CDNS_7246548160514 $T=119630 151025 0 0 $X=119490 $Y=150315
X241 22 VIA1_C_CDNS_7246548160514 $T=125170 118585 0 0 $X=125030 $Y=117875
X242 22 VIA1_C_CDNS_7246548160514 $T=125170 156365 0 0 $X=125030 $Y=155655
X243 2 VIA1_C_CDNS_7246548160514 $T=125870 123925 0 0 $X=125730 $Y=123215
X244 2 VIA1_C_CDNS_7246548160514 $T=125870 151025 0 0 $X=125730 $Y=150315
X245 22 VIA1_C_CDNS_7246548160514 $T=131410 118585 0 0 $X=131270 $Y=117875
X246 22 VIA1_C_CDNS_7246548160514 $T=131410 156365 0 0 $X=131270 $Y=155655
X247 2 VIA1_C_CDNS_7246548160514 $T=132110 123925 0 0 $X=131970 $Y=123215
X248 2 VIA1_C_CDNS_7246548160514 $T=132110 151025 0 0 $X=131970 $Y=150315
X249 22 VIA1_C_CDNS_7246548160514 $T=137650 118585 0 0 $X=137510 $Y=117875
X250 22 VIA1_C_CDNS_7246548160514 $T=137650 156365 0 0 $X=137510 $Y=155655
X251 2 VIA1_C_CDNS_7246548160514 $T=138350 123925 0 0 $X=138210 $Y=123215
X252 2 VIA1_C_CDNS_7246548160514 $T=138350 151025 0 0 $X=138210 $Y=150315
X253 22 VIA1_C_CDNS_7246548160514 $T=143890 118585 0 0 $X=143750 $Y=117875
X254 22 VIA1_C_CDNS_7246548160514 $T=143890 156365 0 0 $X=143750 $Y=155655
X255 2 VIA1_C_CDNS_7246548160514 $T=144590 123925 0 0 $X=144450 $Y=123215
X256 2 VIA1_C_CDNS_7246548160514 $T=144590 151025 0 0 $X=144450 $Y=150315
X257 22 VIA1_C_CDNS_7246548160514 $T=150130 118585 0 0 $X=149990 $Y=117875
X258 22 VIA1_C_CDNS_7246548160514 $T=150130 156365 0 0 $X=149990 $Y=155655
X259 2 VIA1_C_CDNS_7246548160514 $T=150830 123925 0 0 $X=150690 $Y=123215
X260 2 VIA1_C_CDNS_7246548160514 $T=150830 151025 0 0 $X=150690 $Y=150315
X261 18 VIA1_C_CDNS_7246548160514 $T=156370 122145 0 0 $X=156230 $Y=121435
X262 17 VIA1_C_CDNS_7246548160514 $T=156370 152805 0 0 $X=156230 $Y=152095
X263 2 VIA1_C_CDNS_7246548160514 $T=157070 123925 0 0 $X=156930 $Y=123215
X264 2 VIA1_C_CDNS_7246548160514 $T=157070 151025 0 0 $X=156930 $Y=150315
X265 16 VIA1_C_CDNS_7246548160514 $T=162610 116805 0 0 $X=162470 $Y=116095
X266 16 VIA1_C_CDNS_7246548160514 $T=162610 158145 0 0 $X=162470 $Y=157435
X267 2 VIA1_C_CDNS_7246548160514 $T=163310 123925 0 0 $X=163170 $Y=123215
X268 2 VIA1_C_CDNS_7246548160514 $T=163310 151025 0 0 $X=163170 $Y=150315
X269 17 VIA1_C_CDNS_7246548160514 $T=168850 120365 0 0 $X=168710 $Y=119655
X270 18 VIA1_C_CDNS_7246548160514 $T=168850 154585 0 0 $X=168710 $Y=153875
X271 2 VIA1_C_CDNS_7246548160514 $T=169550 123925 0 0 $X=169410 $Y=123215
X272 2 VIA1_C_CDNS_7246548160514 $T=169550 151025 0 0 $X=169410 $Y=150315
X273 22 VIA1_C_CDNS_7246548160514 $T=175090 118585 0 0 $X=174950 $Y=117875
X274 22 VIA1_C_CDNS_7246548160514 $T=175090 156365 0 0 $X=174950 $Y=155655
X275 2 VIA1_C_CDNS_7246548160514 $T=175790 123925 0 0 $X=175650 $Y=123215
X276 2 VIA1_C_CDNS_7246548160514 $T=175790 151025 0 0 $X=175650 $Y=150315
X277 22 VIA1_C_CDNS_7246548160514 $T=181330 118585 0 0 $X=181190 $Y=117875
X278 22 VIA1_C_CDNS_7246548160514 $T=181330 156365 0 0 $X=181190 $Y=155655
X279 2 VIA1_C_CDNS_7246548160514 $T=182030 123925 0 0 $X=181890 $Y=123215
X280 2 VIA1_C_CDNS_7246548160514 $T=182030 151025 0 0 $X=181890 $Y=150315
X281 22 VIA1_C_CDNS_7246548160514 $T=187570 118585 0 0 $X=187430 $Y=117875
X282 22 VIA1_C_CDNS_7246548160514 $T=187570 156365 0 0 $X=187430 $Y=155655
X283 2 VIA1_C_CDNS_7246548160514 $T=188270 123925 0 0 $X=188130 $Y=123215
X284 2 VIA1_C_CDNS_7246548160514 $T=188270 151025 0 0 $X=188130 $Y=150315
X285 22 VIA1_C_CDNS_7246548160514 $T=193810 118585 0 0 $X=193670 $Y=117875
X286 22 VIA1_C_CDNS_7246548160514 $T=193810 156365 0 0 $X=193670 $Y=155655
X287 2 VIA1_C_CDNS_7246548160514 $T=194510 123925 0 0 $X=194370 $Y=123215
X288 2 VIA1_C_CDNS_7246548160514 $T=194510 151025 0 0 $X=194370 $Y=150315
X289 22 VIA1_C_CDNS_7246548160514 $T=200050 118585 0 0 $X=199910 $Y=117875
X290 22 VIA1_C_CDNS_7246548160514 $T=200050 156365 0 0 $X=199910 $Y=155655
X291 2 VIA1_C_CDNS_7246548160514 $T=200750 123925 0 0 $X=200610 $Y=123215
X292 2 VIA1_C_CDNS_7246548160514 $T=200750 151025 0 0 $X=200610 $Y=150315
X293 2 VIA1_C_CDNS_7246548160514 $T=206290 123925 0 0 $X=206150 $Y=123215
X294 2 VIA1_C_CDNS_7246548160514 $T=206290 151025 0 0 $X=206150 $Y=150315
X295 1 VIA1_C_CDNS_7246548160514 $T=231905 19610 0 0 $X=231765 $Y=18900
X296 1 VIA1_C_CDNS_7246548160514 $T=231905 33860 0 0 $X=231765 $Y=33150
X297 20 VIA1_C_CDNS_7246548160514 $T=233445 16050 0 0 $X=233305 $Y=15340
X298 21 VIA1_C_CDNS_7246548160514 $T=233445 35640 0 0 $X=233305 $Y=34930
X299 1 VIA1_C_CDNS_7246548160514 $T=234145 19610 0 0 $X=234005 $Y=18900
X300 1 VIA1_C_CDNS_7246548160514 $T=234145 33860 0 0 $X=234005 $Y=33150
X301 21 VIA1_C_CDNS_7246548160514 $T=235685 17830 0 0 $X=235545 $Y=17120
X302 20 VIA1_C_CDNS_7246548160514 $T=235685 37420 0 0 $X=235545 $Y=36710
X303 24 VIA1_C_CDNS_7246548160515 $T=109005 31610 0 0 $X=108815 $Y=31420
X304 6 VIA1_C_CDNS_7246548160515 $T=109625 32170 0 0 $X=109435 $Y=31980
X305 24 VIA1_C_CDNS_7246548160515 $T=114545 31610 0 0 $X=114355 $Y=31420
X306 6 VIA1_C_CDNS_7246548160515 $T=115165 32170 0 0 $X=114975 $Y=31980
X307 24 VIA1_C_CDNS_7246548160515 $T=120085 31610 0 0 $X=119895 $Y=31420
X308 6 VIA1_C_CDNS_7246548160515 $T=120705 32170 0 0 $X=120515 $Y=31980
X309 24 VIA1_C_CDNS_7246548160515 $T=125625 31610 0 0 $X=125435 $Y=31420
X310 6 VIA1_C_CDNS_7246548160515 $T=126245 32170 0 0 $X=126055 $Y=31980
X311 24 VIA1_C_CDNS_7246548160515 $T=131165 31610 0 0 $X=130975 $Y=31420
X312 6 VIA1_C_CDNS_7246548160515 $T=131785 32170 0 0 $X=131595 $Y=31980
X313 24 VIA1_C_CDNS_7246548160515 $T=136705 31610 0 0 $X=136515 $Y=31420
X314 6 VIA1_C_CDNS_7246548160515 $T=137325 32170 0 0 $X=137135 $Y=31980
X315 24 VIA1_C_CDNS_7246548160515 $T=142245 31610 0 0 $X=142055 $Y=31420
X316 6 VIA1_C_CDNS_7246548160515 $T=142865 32170 0 0 $X=142675 $Y=31980
X317 24 VIA1_C_CDNS_7246548160515 $T=147785 31610 0 0 $X=147595 $Y=31420
X318 6 VIA1_C_CDNS_7246548160515 $T=148405 32170 0 0 $X=148215 $Y=31980
X319 24 VIA1_C_CDNS_7246548160515 $T=153325 31610 0 0 $X=153135 $Y=31420
X320 6 VIA1_C_CDNS_7246548160515 $T=153945 32170 0 0 $X=153755 $Y=31980
X321 24 VIA1_C_CDNS_7246548160515 $T=163595 31610 0 0 $X=163405 $Y=31420
X322 6 VIA1_C_CDNS_7246548160515 $T=164105 32170 0 0 $X=163915 $Y=31980
X323 24 VIA1_C_CDNS_7246548160515 $T=169135 31610 0 0 $X=168945 $Y=31420
X324 6 VIA1_C_CDNS_7246548160515 $T=169645 32170 0 0 $X=169455 $Y=31980
X325 24 VIA1_C_CDNS_7246548160515 $T=174675 31610 0 0 $X=174485 $Y=31420
X326 6 VIA1_C_CDNS_7246548160515 $T=175185 32170 0 0 $X=174995 $Y=31980
X327 24 VIA1_C_CDNS_7246548160515 $T=180215 31610 0 0 $X=180025 $Y=31420
X328 6 VIA1_C_CDNS_7246548160515 $T=180725 32170 0 0 $X=180535 $Y=31980
X329 24 VIA1_C_CDNS_7246548160515 $T=185755 31610 0 0 $X=185565 $Y=31420
X330 6 VIA1_C_CDNS_7246548160515 $T=186265 32170 0 0 $X=186075 $Y=31980
X331 24 VIA1_C_CDNS_7246548160515 $T=191295 31610 0 0 $X=191105 $Y=31420
X332 6 VIA1_C_CDNS_7246548160515 $T=191805 32170 0 0 $X=191615 $Y=31980
X333 24 VIA1_C_CDNS_7246548160515 $T=196835 31610 0 0 $X=196645 $Y=31420
X334 6 VIA1_C_CDNS_7246548160515 $T=197345 32170 0 0 $X=197155 $Y=31980
X335 24 VIA1_C_CDNS_7246548160515 $T=202375 31610 0 0 $X=202185 $Y=31420
X336 6 VIA1_C_CDNS_7246548160515 $T=202885 32170 0 0 $X=202695 $Y=31980
X337 24 VIA1_C_CDNS_7246548160515 $T=207915 31610 0 0 $X=207725 $Y=31420
X338 6 VIA1_C_CDNS_7246548160515 $T=208425 32170 0 0 $X=208235 $Y=31980
X339 17 1 ND_C_CDNS_7246548160516 $T=131350 17825 0 0 $X=106195 $Y=17420
X340 18 1 ND_C_CDNS_7246548160516 $T=131350 45950 0 0 $X=106195 $Y=45545
X341 18 1 ND_C_CDNS_7246548160516 $T=185880 16050 0 0 $X=160725 $Y=15645
X342 17 1 ND_C_CDNS_7246548160516 $T=185880 47720 0 0 $X=160725 $Y=47315
X343 1 VIA2_C_CDNS_7246548160517 $T=112085 14270 0 0 $X=111685 $Y=13560
X344 1 VIA2_C_CDNS_7246548160517 $T=112085 49510 0 0 $X=111685 $Y=48800
X345 1 VIA2_C_CDNS_7246548160517 $T=123165 14270 0 0 $X=122765 $Y=13560
X346 1 VIA2_C_CDNS_7246548160517 $T=123165 49510 0 0 $X=122765 $Y=48800
X347 1 VIA2_C_CDNS_7246548160517 $T=134245 14270 0 0 $X=133845 $Y=13560
X348 1 VIA2_C_CDNS_7246548160517 $T=134245 49510 0 0 $X=133845 $Y=48800
X349 1 VIA2_C_CDNS_7246548160517 $T=145325 14270 0 0 $X=144925 $Y=13560
X350 1 VIA2_C_CDNS_7246548160517 $T=145325 49510 0 0 $X=144925 $Y=48800
X351 1 VIA2_C_CDNS_7246548160517 $T=156405 14270 0 0 $X=156005 $Y=13560
X352 1 VIA2_C_CDNS_7246548160517 $T=156405 49510 0 0 $X=156005 $Y=48800
X353 1 VIA2_C_CDNS_7246548160517 $T=166365 14270 0 0 $X=165965 $Y=13560
X354 1 VIA2_C_CDNS_7246548160517 $T=166365 49510 0 0 $X=165965 $Y=48800
X355 1 VIA2_C_CDNS_7246548160517 $T=177445 14270 0 0 $X=177045 $Y=13560
X356 1 VIA2_C_CDNS_7246548160517 $T=177445 49510 0 0 $X=177045 $Y=48800
X357 1 VIA2_C_CDNS_7246548160517 $T=188525 14270 0 0 $X=188125 $Y=13560
X358 1 VIA2_C_CDNS_7246548160517 $T=188525 49510 0 0 $X=188125 $Y=48800
X359 1 VIA2_C_CDNS_7246548160517 $T=199605 14270 0 0 $X=199205 $Y=13560
X360 1 VIA2_C_CDNS_7246548160517 $T=199605 49510 0 0 $X=199205 $Y=48800
X361 1 VIA2_C_CDNS_7246548160517 $T=210685 14270 0 0 $X=210285 $Y=13560
X362 1 VIA2_C_CDNS_7246548160517 $T=210685 49510 0 0 $X=210285 $Y=48800
X363 3 VIA1_C_CDNS_7246548160518 $T=13505 83830 0 0 $X=13015 $Y=83600
X364 3 VIA1_C_CDNS_7246548160518 $T=13505 86055 0 0 $X=13015 $Y=85825
X365 5 VIA1_C_CDNS_7246548160518 $T=17705 83830 0 0 $X=17215 $Y=83600
X366 5 VIA1_C_CDNS_7246548160518 $T=17705 86055 0 0 $X=17215 $Y=85825
X367 25 VIA1_C_CDNS_7246548160519 $T=23615 88310 0 0 $X=22865 $Y=88080
X368 26 VIA1_C_CDNS_7246548160519 $T=24350 86955 0 0 $X=23600 $Y=86725
X369 1 VIA1_C_CDNS_7246548160521 $T=105815 12260 0 0 $X=103025 $Y=11060
X370 1 VIA1_C_CDNS_7246548160521 $T=211445 12030 0 0 $X=208655 $Y=10830
X371 1 VIA2_C_CDNS_7246548160522 $T=105815 12260 0 0 $X=103025 $Y=11060
X372 1 VIA2_C_CDNS_7246548160522 $T=211445 12030 0 0 $X=208655 $Y=10830
X373 17 VIA1_C_CDNS_7246548160523 $T=101790 44390 0 0 $X=101040 $Y=42080
X374 18 VIA1_C_CDNS_7246548160523 $T=215715 44390 0 0 $X=214965 $Y=42080
X375 1 VIA1_C_CDNS_7246548160524 $T=243980 19610 0 0 $X=241930 $Y=18860
X376 23 VIA1_C_CDNS_7246548160524 $T=311195 26360 0 0 $X=309145 $Y=25610
X377 9 VIA1_C_CDNS_7246548160524 $T=315635 26360 0 0 $X=313585 $Y=25610
X378 23 VIA1_C_CDNS_7246548160524 $T=324920 82035 0 0 $X=322870 $Y=81285
X379 19 VIA2_C_CDNS_7246548160525 $T=92185 100410 0 0 $X=89615 $Y=99660
X380 19 VIA2_C_CDNS_7246548160525 $T=249890 17585 0 0 $X=247320 $Y=16835
X381 2 1 VIA2_C_CDNS_7246548160527 $T=110885 161700 0 0 $X=108315 $Y=160170
X382 2 1 VIA2_C_CDNS_7246548160527 $T=208825 161700 0 0 $X=206255 $Y=160170
X383 2 1 VIA1_C_CDNS_7246548160528 $T=105735 160860 0 0 $X=97965 $Y=160110
X384 2 1 VIA1_C_CDNS_7246548160528 $T=213285 160860 0 0 $X=205515 $Y=160110
X385 27 VIA2_C_CDNS_7246548160535 $T=259810 122590 0 0 $X=259320 $Y=120540
X386 27 VIA1_C_CDNS_7246548160536 $T=259810 122590 0 0 $X=259320 $Y=120540
X387 23 VIA3_C_CDNS_7246548160537 $T=311195 26360 0 0 $X=309145 $Y=25610
X388 9 VIA3_C_CDNS_7246548160537 $T=315635 26360 0 0 $X=313585 $Y=25610
X389 23 VIA3_C_CDNS_7246548160537 $T=324920 82035 0 0 $X=322870 $Y=81285
X390 10 VIA1_C_CDNS_7246548160539 $T=354705 81715 0 0 $X=352655 $Y=81225
X391 19 VIA2_C_CDNS_7246548160541 $T=259880 101230 0 0 $X=259650 $Y=99180
X392 6 VIA2_C_CDNS_7246548160543 $T=98240 32160 0 0 $X=97490 $Y=31410
X393 19 VIA2_C_CDNS_7246548160543 $T=259885 73765 0 0 $X=259135 $Y=73015
X394 7 VIATP_C_CDNS_7246548160545 $T=376900 51365 0 0 $X=376110 $Y=50835
X395 7 VIATP_C_CDNS_7246548160545 $T=376900 147425 0 0 $X=376110 $Y=146895
X396 11 VIATP_C_CDNS_7246548160545 $T=557055 51365 0 0 $X=556265 $Y=50835
X397 11 VIATP_C_CDNS_7246548160545 $T=557055 147425 0 0 $X=556265 $Y=146895
X398 7 VIATP_C_CDNS_7246548160549 $T=433355 51365 0 0 $X=432695 $Y=50835
X399 7 VIATP_C_CDNS_7246548160549 $T=433355 147425 0 0 $X=432695 $Y=146895
X400 11 VIATP_C_CDNS_7246548160549 $T=500600 51365 0 0 $X=499940 $Y=50835
X401 11 VIATP_C_CDNS_7246548160549 $T=500600 147425 0 0 $X=499940 $Y=146895
X402 3 VIA2_C_CDNS_7246548160557 $T=13245 83830 0 0 $X=12495 $Y=83600
X403 5 VIA2_C_CDNS_7246548160557 $T=17445 83830 0 0 $X=16695 $Y=83600
X404 1 20 19 ne3_CDNS_724654816050 $T=248120 21400 0 0 $X=247320 $Y=21000
X405 8 23 9 19 nedia_CDNS_724654816051 $T=282450 37820 0 0 $X=266230 $Y=18430
X406 1 26 12 ne3_CDNS_724654816052 $T=25060 81535 0 0 $X=24260 $Y=80955
X407 1 25 20 ne3_CDNS_724654816052 $T=30635 81535 0 0 $X=29835 $Y=80955
X408 23 9 8 rpp1k1_3_CDNS_724654816053 $T=317545 27490 0 90 $X=309065 $Y=26550
X409 8 11 7 23 nedia_CDNS_724654816054 $T=441980 141045 0 270 $X=422590 $Y=41525
X410 12 4 4 1 ne3_CDNS_724654816055 $T=8060 64240 0 0 $X=7260 $Y=63840
X411 13 4 14 1 ne3_CDNS_724654816055 $T=33845 64240 0 0 $X=33045 $Y=63840
X412 15 4 16 1 ne3_CDNS_724654816055 $T=59570 64240 0 0 $X=58770 $Y=63840
X413 2 14 19 2 1 pe3_CDNS_724654816056 $T=63965 94930 0 180 $X=61455 $Y=83900
X414 2 14 19 2 1 pe3_CDNS_724654816056 $T=66205 94930 0 180 $X=63695 $Y=83900
X415 2 14 14 2 1 pe3_CDNS_724654816056 $T=68445 94930 0 180 $X=65935 $Y=83900
X416 2 14 19 2 1 pe3_CDNS_724654816056 $T=70685 94930 0 180 $X=68175 $Y=83900
X417 2 14 19 2 1 pe3_CDNS_724654816056 $T=72925 94930 0 180 $X=70415 $Y=83900
X418 2 3 26 1 pe3_CDNS_724654816057 $T=15530 89865 0 180 $X=13480 $Y=86295
X419 2 5 25 1 pe3_CDNS_724654816057 $T=19690 89865 0 180 $X=17640 $Y=86295
X420 9 11 8 rpp1k1_3_CDNS_724654816058 $T=558265 45130 0 90 $X=515365 $Y=41970
X421 2 2 2 2 1 pe3_CDNS_7246548160511 $T=109700 69700 0 0 $X=108190 $Y=68670
X422 2 2 2 2 1 pe3_CDNS_7246548160511 $T=109700 93320 1 0 $X=108190 $Y=82290
X423 2 2 2 2 1 pe3_CDNS_7246548160511 $T=113660 125985 0 0 $X=112150 $Y=124955
X424 2 2 2 2 1 pe3_CDNS_7246548160511 $T=113660 148965 1 0 $X=112150 $Y=137935
X425 22 18 20 2 1 pe3_CDNS_7246548160511 $T=115940 69700 0 0 $X=114430 $Y=68670
X426 22 17 21 2 1 pe3_CDNS_7246548160511 $T=115940 93320 1 0 $X=114430 $Y=82290
X427 2 16 22 2 1 pe3_CDNS_7246548160511 $T=119900 125985 0 0 $X=118390 $Y=124955
X428 2 16 22 2 1 pe3_CDNS_7246548160511 $T=119900 148965 1 0 $X=118390 $Y=137935
X429 22 17 21 2 1 pe3_CDNS_7246548160511 $T=122180 69700 0 0 $X=120670 $Y=68670
X430 22 18 20 2 1 pe3_CDNS_7246548160511 $T=122180 93320 1 0 $X=120670 $Y=82290
X431 2 16 22 2 1 pe3_CDNS_7246548160511 $T=126140 125985 0 0 $X=124630 $Y=124955
X432 2 16 22 2 1 pe3_CDNS_7246548160511 $T=126140 148965 1 0 $X=124630 $Y=137935
X433 22 18 20 2 1 pe3_CDNS_7246548160511 $T=128420 69700 0 0 $X=126910 $Y=68670
X434 22 17 21 2 1 pe3_CDNS_7246548160511 $T=128420 93320 1 0 $X=126910 $Y=82290
X435 2 16 22 2 1 pe3_CDNS_7246548160511 $T=132380 125985 0 0 $X=130870 $Y=124955
X436 2 16 22 2 1 pe3_CDNS_7246548160511 $T=132380 148965 1 0 $X=130870 $Y=137935
X437 22 17 21 2 1 pe3_CDNS_7246548160511 $T=134660 69700 0 0 $X=133150 $Y=68670
X438 22 18 20 2 1 pe3_CDNS_7246548160511 $T=134660 93320 1 0 $X=133150 $Y=82290
X439 2 16 22 2 1 pe3_CDNS_7246548160511 $T=138620 125985 0 0 $X=137110 $Y=124955
X440 2 16 22 2 1 pe3_CDNS_7246548160511 $T=138620 148965 1 0 $X=137110 $Y=137935
X441 22 18 20 2 1 pe3_CDNS_7246548160511 $T=140900 69700 0 0 $X=139390 $Y=68670
X442 22 17 21 2 1 pe3_CDNS_7246548160511 $T=140900 93320 1 0 $X=139390 $Y=82290
X443 2 16 22 2 1 pe3_CDNS_7246548160511 $T=144860 125985 0 0 $X=143350 $Y=124955
X444 2 16 22 2 1 pe3_CDNS_7246548160511 $T=144860 148965 1 0 $X=143350 $Y=137935
X445 22 17 21 2 1 pe3_CDNS_7246548160511 $T=147140 69700 0 0 $X=145630 $Y=68670
X446 22 18 20 2 1 pe3_CDNS_7246548160511 $T=147140 93320 1 0 $X=145630 $Y=82290
X447 2 16 18 2 1 pe3_CDNS_7246548160511 $T=151100 125985 0 0 $X=149590 $Y=124955
X448 2 16 17 2 1 pe3_CDNS_7246548160511 $T=151100 148965 1 0 $X=149590 $Y=137935
X449 22 18 20 2 1 pe3_CDNS_7246548160511 $T=153380 69700 0 0 $X=151870 $Y=68670
X450 22 17 21 2 1 pe3_CDNS_7246548160511 $T=153380 93320 1 0 $X=151870 $Y=82290
X451 2 16 16 2 1 pe3_CDNS_7246548160511 $T=157340 125985 0 0 $X=155830 $Y=124955
X452 2 16 16 2 1 pe3_CDNS_7246548160511 $T=157340 148965 1 0 $X=155830 $Y=137935
X453 22 17 21 2 1 pe3_CDNS_7246548160511 $T=159620 69700 0 0 $X=158110 $Y=68670
X454 22 18 20 2 1 pe3_CDNS_7246548160511 $T=159620 93320 1 0 $X=158110 $Y=82290
X455 2 16 17 2 1 pe3_CDNS_7246548160511 $T=163580 125985 0 0 $X=162070 $Y=124955
X456 2 16 18 2 1 pe3_CDNS_7246548160511 $T=163580 148965 1 0 $X=162070 $Y=137935
X457 22 18 20 2 1 pe3_CDNS_7246548160511 $T=165860 69700 0 0 $X=164350 $Y=68670
X458 22 17 21 2 1 pe3_CDNS_7246548160511 $T=165860 93320 1 0 $X=164350 $Y=82290
X459 2 16 22 2 1 pe3_CDNS_7246548160511 $T=169820 125985 0 0 $X=168310 $Y=124955
X460 2 16 22 2 1 pe3_CDNS_7246548160511 $T=169820 148965 1 0 $X=168310 $Y=137935
X461 22 17 21 2 1 pe3_CDNS_7246548160511 $T=172100 69700 0 0 $X=170590 $Y=68670
X462 22 18 20 2 1 pe3_CDNS_7246548160511 $T=172100 93320 1 0 $X=170590 $Y=82290
X463 2 16 22 2 1 pe3_CDNS_7246548160511 $T=176060 125985 0 0 $X=174550 $Y=124955
X464 2 16 22 2 1 pe3_CDNS_7246548160511 $T=176060 148965 1 0 $X=174550 $Y=137935
X465 22 18 20 2 1 pe3_CDNS_7246548160511 $T=178340 69700 0 0 $X=176830 $Y=68670
X466 22 17 21 2 1 pe3_CDNS_7246548160511 $T=178340 93320 1 0 $X=176830 $Y=82290
X467 2 16 22 2 1 pe3_CDNS_7246548160511 $T=182300 125985 0 0 $X=180790 $Y=124955
X468 2 16 22 2 1 pe3_CDNS_7246548160511 $T=182300 148965 1 0 $X=180790 $Y=137935
X469 22 17 21 2 1 pe3_CDNS_7246548160511 $T=184580 69700 0 0 $X=183070 $Y=68670
X470 22 18 20 2 1 pe3_CDNS_7246548160511 $T=184580 93320 1 0 $X=183070 $Y=82290
X471 2 16 22 2 1 pe3_CDNS_7246548160511 $T=188540 125985 0 0 $X=187030 $Y=124955
X472 2 16 22 2 1 pe3_CDNS_7246548160511 $T=188540 148965 1 0 $X=187030 $Y=137935
X473 22 18 20 2 1 pe3_CDNS_7246548160511 $T=190820 69700 0 0 $X=189310 $Y=68670
X474 22 17 21 2 1 pe3_CDNS_7246548160511 $T=190820 93320 1 0 $X=189310 $Y=82290
X475 2 16 22 2 1 pe3_CDNS_7246548160511 $T=194780 125985 0 0 $X=193270 $Y=124955
X476 2 16 22 2 1 pe3_CDNS_7246548160511 $T=194780 148965 1 0 $X=193270 $Y=137935
X477 22 17 21 2 1 pe3_CDNS_7246548160511 $T=197060 69700 0 0 $X=195550 $Y=68670
X478 22 18 20 2 1 pe3_CDNS_7246548160511 $T=197060 93320 1 0 $X=195550 $Y=82290
X479 2 2 2 2 1 pe3_CDNS_7246548160511 $T=201020 125985 0 0 $X=199510 $Y=124955
X480 2 2 2 2 1 pe3_CDNS_7246548160511 $T=201020 148965 1 0 $X=199510 $Y=137935
X481 2 2 2 2 1 pe3_CDNS_7246548160511 $T=203300 69700 0 0 $X=201790 $Y=68670
X482 2 2 2 2 1 pe3_CDNS_7246548160511 $T=203300 93320 1 0 $X=201790 $Y=82290
X483 1 1 1 ne3_CDNS_7246548160512 $T=17420 20740 0 0 $X=16620 $Y=20340
X484 1 1 1 ne3_CDNS_7246548160512 $T=17420 42860 1 0 $X=16620 $Y=32290
X485 1 12 15 ne3_CDNS_7246548160512 $T=28660 20740 0 0 $X=27860 $Y=20340
X486 1 12 15 ne3_CDNS_7246548160512 $T=28660 42860 1 0 $X=27860 $Y=32290
X487 1 12 12 ne3_CDNS_7246548160512 $T=39900 20740 0 0 $X=39100 $Y=20340
X488 1 12 12 ne3_CDNS_7246548160512 $T=39900 42860 1 0 $X=39100 $Y=32290
X489 1 12 13 ne3_CDNS_7246548160512 $T=51140 20740 0 0 $X=50340 $Y=20340
X490 1 12 13 ne3_CDNS_7246548160512 $T=51140 42860 1 0 $X=50340 $Y=32290
X491 1 1 1 ne3_CDNS_7246548160512 $T=62380 20740 0 0 $X=61580 $Y=20340
X492 1 1 1 ne3_CDNS_7246548160512 $T=62380 42860 1 0 $X=61580 $Y=32290
X493 1 21 20 ne3_CDNS_7246548160513 $T=232175 21040 0 0 $X=231375 $Y=20640
X494 1 21 21 ne3_CDNS_7246548160513 $T=232175 32430 1 0 $X=231375 $Y=26860
X495 1 21 21 ne3_CDNS_7246548160513 $T=234415 21040 0 0 $X=233615 $Y=20640
X496 1 21 20 ne3_CDNS_7246548160513 $T=234415 32430 1 0 $X=233615 $Y=26860
X497 17 6 1 pe3_CDNS_7246548160514 $T=106815 19890 0 0 $X=105305 $Y=18860
X498 18 24 1 pe3_CDNS_7246548160514 $T=106815 43890 1 0 $X=105305 $Y=32860
X499 18 24 1 pe3_CDNS_7246548160514 $T=161095 19890 0 0 $X=159585 $Y=18860
X500 17 6 1 pe3_CDNS_7246548160514 $T=161095 43890 1 0 $X=159585 $Y=32860
X501 7 24 1 rpp1k1_3_CDNS_7246548160515 $T=229190 61300 0 90 $X=226970 $Y=60360
X502 7 24 1 rpp1k1_3_CDNS_7246548160515 $T=232060 61300 0 90 $X=229840 $Y=60360
X503 7 24 1 rpp1k1_3_CDNS_7246548160515 $T=234930 61300 0 90 $X=232710 $Y=60360
X504 7 24 1 rpp1k1_3_CDNS_7246548160515 $T=237800 61300 0 90 $X=235580 $Y=60360
X505 7 24 1 rpp1k1_3_CDNS_7246548160515 $T=240670 61300 0 90 $X=238450 $Y=60360
X506 7 24 1 rpp1k1_3_CDNS_7246548160515 $T=243540 61300 0 90 $X=241320 $Y=60360
X507 7 24 1 rpp1k1_3_CDNS_7246548160515 $T=246410 61300 0 90 $X=244190 $Y=60360
X508 7 24 1 rpp1k1_3_CDNS_7246548160515 $T=249280 61300 0 90 $X=247060 $Y=60360
X509 7 24 1 rpp1k1_3_CDNS_7246548160515 $T=252150 61300 0 90 $X=249930 $Y=60360
X510 19 27 2 1 rpp1k1_3_CDNS_7246548160516 $T=255085 124550 0 180 $X=228430 $Y=99030
X511 10 23 8 rpp1k1_3_CDNS_7246548160517 $T=322885 76685 0 270 $X=322665 $Y=25845
X512 1 3 26 ne3_CDNS_7246548160518 $T=14340 81020 0 0 $X=13540 $Y=80620
X513 1 5 25 ne3_CDNS_7246548160518 $T=18500 81020 0 0 $X=17700 $Y=80620
X514 7 MASCO__X1 $T=432695 51895 0 0 $X=432695 $Y=51895
X515 7 MASCO__X1 $T=432695 56895 0 0 $X=432695 $Y=56895
X516 7 MASCO__X1 $T=432695 61895 0 0 $X=432695 $Y=61895
X517 7 MASCO__X1 $T=432695 66895 0 0 $X=432695 $Y=66895
X518 7 MASCO__X1 $T=432695 71895 0 0 $X=432695 $Y=71895
X519 7 MASCO__X1 $T=432695 76895 0 0 $X=432695 $Y=76895
X520 7 MASCO__X1 $T=432695 81895 0 0 $X=432695 $Y=81895
X521 7 MASCO__X1 $T=432695 86895 0 0 $X=432695 $Y=86895
X522 7 MASCO__X1 $T=432695 91895 0 0 $X=432695 $Y=91895
X523 7 MASCO__X1 $T=432695 96895 0 0 $X=432695 $Y=96895
X524 7 MASCO__X1 $T=432695 101895 0 0 $X=432695 $Y=101895
X525 7 MASCO__X1 $T=432695 106895 0 0 $X=432695 $Y=106895
X526 7 MASCO__X1 $T=432695 111895 0 0 $X=432695 $Y=111895
X527 7 MASCO__X1 $T=432695 116895 0 0 $X=432695 $Y=116895
X528 7 MASCO__X1 $T=432695 121895 0 0 $X=432695 $Y=121895
X529 7 MASCO__X1 $T=432695 126895 0 0 $X=432695 $Y=126895
X530 7 MASCO__X1 $T=432695 131895 0 0 $X=432695 $Y=131895
X531 7 MASCO__X1 $T=432695 136895 0 0 $X=432695 $Y=136895
X532 7 MASCO__X1 $T=432695 141895 0 0 $X=432695 $Y=141895
X533 11 MASCO__X1 $T=499940 51895 0 0 $X=499940 $Y=51895
X534 11 MASCO__X1 $T=499940 56895 0 0 $X=499940 $Y=56895
X535 11 MASCO__X1 $T=499940 61895 0 0 $X=499940 $Y=61895
X536 11 MASCO__X1 $T=499940 66895 0 0 $X=499940 $Y=66895
X537 11 MASCO__X1 $T=499940 71895 0 0 $X=499940 $Y=71895
X538 11 MASCO__X1 $T=499940 76895 0 0 $X=499940 $Y=76895
X539 11 MASCO__X1 $T=499940 81895 0 0 $X=499940 $Y=81895
X540 11 MASCO__X1 $T=499940 86895 0 0 $X=499940 $Y=86895
X541 11 MASCO__X1 $T=499940 91895 0 0 $X=499940 $Y=91895
X542 11 MASCO__X1 $T=499940 96895 0 0 $X=499940 $Y=96895
X543 11 MASCO__X1 $T=499940 101895 0 0 $X=499940 $Y=101895
X544 11 MASCO__X1 $T=499940 106895 0 0 $X=499940 $Y=106895
X545 11 MASCO__X1 $T=499940 111895 0 0 $X=499940 $Y=111895
X546 11 MASCO__X1 $T=499940 116895 0 0 $X=499940 $Y=116895
X547 11 MASCO__X1 $T=499940 121895 0 0 $X=499940 $Y=121895
X548 11 MASCO__X1 $T=499940 126895 0 0 $X=499940 $Y=126895
X549 11 MASCO__X1 $T=499940 131895 0 0 $X=499940 $Y=131895
X550 11 MASCO__X1 $T=499940 136895 0 0 $X=499940 $Y=136895
X551 11 MASCO__X1 $T=499940 141895 0 0 $X=499940 $Y=141895
X552 7 MASCO__X2 $T=376110 51895 0 0 $X=376110 $Y=51895
X553 7 MASCO__X2 $T=376110 56895 0 0 $X=376110 $Y=56895
X554 7 MASCO__X2 $T=376110 61895 0 0 $X=376110 $Y=61895
X555 7 MASCO__X2 $T=376110 66895 0 0 $X=376110 $Y=66895
X556 7 MASCO__X2 $T=376110 71895 0 0 $X=376110 $Y=71895
X557 7 MASCO__X2 $T=376110 76895 0 0 $X=376110 $Y=76895
X558 7 MASCO__X2 $T=376110 81895 0 0 $X=376110 $Y=81895
X559 7 MASCO__X2 $T=376110 86895 0 0 $X=376110 $Y=86895
X560 7 MASCO__X2 $T=376110 91895 0 0 $X=376110 $Y=91895
X561 7 MASCO__X2 $T=376110 96895 0 0 $X=376110 $Y=96895
X562 7 MASCO__X2 $T=376110 101895 0 0 $X=376110 $Y=101895
X563 7 MASCO__X2 $T=376110 106895 0 0 $X=376110 $Y=106895
X564 7 MASCO__X2 $T=376110 111895 0 0 $X=376110 $Y=111895
X565 7 MASCO__X2 $T=376110 116895 0 0 $X=376110 $Y=116895
X566 7 MASCO__X2 $T=376110 121895 0 0 $X=376110 $Y=121895
X567 7 MASCO__X2 $T=376110 126895 0 0 $X=376110 $Y=126895
X568 7 MASCO__X2 $T=376110 131895 0 0 $X=376110 $Y=131895
X569 7 MASCO__X2 $T=376110 136895 0 0 $X=376110 $Y=136895
X570 7 MASCO__X2 $T=376110 141895 0 0 $X=376110 $Y=141895
X571 11 MASCO__X2 $T=556265 51895 0 0 $X=556265 $Y=51895
X572 11 MASCO__X2 $T=556265 56895 0 0 $X=556265 $Y=56895
X573 11 MASCO__X2 $T=556265 61895 0 0 $X=556265 $Y=61895
X574 11 MASCO__X2 $T=556265 66895 0 0 $X=556265 $Y=66895
X575 11 MASCO__X2 $T=556265 71895 0 0 $X=556265 $Y=71895
X576 11 MASCO__X2 $T=556265 76895 0 0 $X=556265 $Y=76895
X577 11 MASCO__X2 $T=556265 81895 0 0 $X=556265 $Y=81895
X578 11 MASCO__X2 $T=556265 86895 0 0 $X=556265 $Y=86895
X579 11 MASCO__X2 $T=556265 91895 0 0 $X=556265 $Y=91895
X580 11 MASCO__X2 $T=556265 96895 0 0 $X=556265 $Y=96895
X581 11 MASCO__X2 $T=556265 101895 0 0 $X=556265 $Y=101895
X582 11 MASCO__X2 $T=556265 106895 0 0 $X=556265 $Y=106895
X583 11 MASCO__X2 $T=556265 111895 0 0 $X=556265 $Y=111895
X584 11 MASCO__X2 $T=556265 116895 0 0 $X=556265 $Y=116895
X585 11 MASCO__X2 $T=556265 121895 0 0 $X=556265 $Y=121895
X586 11 MASCO__X2 $T=556265 126895 0 0 $X=556265 $Y=126895
X587 11 MASCO__X2 $T=556265 131895 0 0 $X=556265 $Y=131895
X588 11 MASCO__X2 $T=556265 136895 0 0 $X=556265 $Y=136895
X589 11 MASCO__X2 $T=556265 141895 0 0 $X=556265 $Y=141895
X590 7 MASCO__Y6 $T=378695 51895 0 0 $X=378695 $Y=51895
X591 7 MASCO__Y6 $T=378695 56895 0 0 $X=378695 $Y=56895
X592 7 MASCO__Y6 $T=378695 61895 0 0 $X=378695 $Y=61895
X593 7 MASCO__Y6 $T=378695 66895 0 0 $X=378695 $Y=66895
X594 7 MASCO__Y6 $T=378695 71895 0 0 $X=378695 $Y=71895
X595 7 MASCO__Y6 $T=378695 76895 0 0 $X=378695 $Y=76895
X596 7 MASCO__Y6 $T=378695 81895 0 0 $X=378695 $Y=81895
X597 7 MASCO__Y6 $T=378695 86895 0 0 $X=378695 $Y=86895
X598 7 MASCO__Y6 $T=378695 91895 0 0 $X=378695 $Y=91895
X599 7 MASCO__Y6 $T=378695 96895 0 0 $X=378695 $Y=96895
X600 7 MASCO__Y6 $T=378695 101895 0 0 $X=378695 $Y=101895
X601 7 MASCO__Y6 $T=378695 106895 0 0 $X=378695 $Y=106895
X602 7 MASCO__Y6 $T=378695 111895 0 0 $X=378695 $Y=111895
X603 7 MASCO__Y6 $T=378695 116895 0 0 $X=378695 $Y=116895
X604 7 MASCO__Y6 $T=378695 121895 0 0 $X=378695 $Y=121895
X605 7 MASCO__Y6 $T=378695 126895 0 0 $X=378695 $Y=126895
X606 7 MASCO__Y6 $T=378695 131895 0 0 $X=378695 $Y=131895
X607 7 MASCO__Y6 $T=378695 136895 0 0 $X=378695 $Y=136895
X608 7 MASCO__Y6 $T=378695 141895 0 0 $X=378695 $Y=141895
X609 7 MASCO__Y6 $T=396695 51895 0 0 $X=396695 $Y=51895
X610 7 MASCO__Y6 $T=396695 56895 0 0 $X=396695 $Y=56895
X611 7 MASCO__Y6 $T=396695 61895 0 0 $X=396695 $Y=61895
X612 7 MASCO__Y6 $T=396695 66895 0 0 $X=396695 $Y=66895
X613 7 MASCO__Y6 $T=396695 71895 0 0 $X=396695 $Y=71895
X614 7 MASCO__Y6 $T=396695 76895 0 0 $X=396695 $Y=76895
X615 7 MASCO__Y6 $T=396695 81895 0 0 $X=396695 $Y=81895
X616 7 MASCO__Y6 $T=396695 86895 0 0 $X=396695 $Y=86895
X617 7 MASCO__Y6 $T=396695 91895 0 0 $X=396695 $Y=91895
X618 7 MASCO__Y6 $T=396695 96895 0 0 $X=396695 $Y=96895
X619 7 MASCO__Y6 $T=396695 101895 0 0 $X=396695 $Y=101895
X620 7 MASCO__Y6 $T=396695 106895 0 0 $X=396695 $Y=106895
X621 7 MASCO__Y6 $T=396695 111895 0 0 $X=396695 $Y=111895
X622 7 MASCO__Y6 $T=396695 116895 0 0 $X=396695 $Y=116895
X623 7 MASCO__Y6 $T=396695 121895 0 0 $X=396695 $Y=121895
X624 7 MASCO__Y6 $T=396695 126895 0 0 $X=396695 $Y=126895
X625 7 MASCO__Y6 $T=396695 131895 0 0 $X=396695 $Y=131895
X626 7 MASCO__Y6 $T=396695 136895 0 0 $X=396695 $Y=136895
X627 7 MASCO__Y6 $T=396695 141895 0 0 $X=396695 $Y=141895
X628 7 MASCO__Y6 $T=414695 51895 0 0 $X=414695 $Y=51895
X629 7 MASCO__Y6 $T=414695 56895 0 0 $X=414695 $Y=56895
X630 7 MASCO__Y6 $T=414695 61895 0 0 $X=414695 $Y=61895
X631 7 MASCO__Y6 $T=414695 66895 0 0 $X=414695 $Y=66895
X632 7 MASCO__Y6 $T=414695 71895 0 0 $X=414695 $Y=71895
X633 7 MASCO__Y6 $T=414695 76895 0 0 $X=414695 $Y=76895
X634 7 MASCO__Y6 $T=414695 81895 0 0 $X=414695 $Y=81895
X635 7 MASCO__Y6 $T=414695 86895 0 0 $X=414695 $Y=86895
X636 7 MASCO__Y6 $T=414695 91895 0 0 $X=414695 $Y=91895
X637 7 MASCO__Y6 $T=414695 96895 0 0 $X=414695 $Y=96895
X638 7 MASCO__Y6 $T=414695 101895 0 0 $X=414695 $Y=101895
X639 7 MASCO__Y6 $T=414695 106895 0 0 $X=414695 $Y=106895
X640 7 MASCO__Y6 $T=414695 111895 0 0 $X=414695 $Y=111895
X641 7 MASCO__Y6 $T=414695 116895 0 0 $X=414695 $Y=116895
X642 7 MASCO__Y6 $T=414695 121895 0 0 $X=414695 $Y=121895
X643 7 MASCO__Y6 $T=414695 126895 0 0 $X=414695 $Y=126895
X644 7 MASCO__Y6 $T=414695 131895 0 0 $X=414695 $Y=131895
X645 7 MASCO__Y6 $T=414695 136895 0 0 $X=414695 $Y=136895
X646 7 MASCO__Y6 $T=414695 141895 0 0 $X=414695 $Y=141895
X647 11 MASCO__Y6 $T=502265 51895 0 0 $X=502265 $Y=51895
X648 11 MASCO__Y6 $T=502265 56895 0 0 $X=502265 $Y=56895
X649 11 MASCO__Y6 $T=502265 61895 0 0 $X=502265 $Y=61895
X650 11 MASCO__Y6 $T=502265 66895 0 0 $X=502265 $Y=66895
X651 11 MASCO__Y6 $T=502265 71895 0 0 $X=502265 $Y=71895
X652 11 MASCO__Y6 $T=502265 76895 0 0 $X=502265 $Y=76895
X653 11 MASCO__Y6 $T=502265 81895 0 0 $X=502265 $Y=81895
X654 11 MASCO__Y6 $T=502265 86895 0 0 $X=502265 $Y=86895
X655 11 MASCO__Y6 $T=502265 91895 0 0 $X=502265 $Y=91895
X656 11 MASCO__Y6 $T=502265 96895 0 0 $X=502265 $Y=96895
X657 11 MASCO__Y6 $T=502265 101895 0 0 $X=502265 $Y=101895
X658 11 MASCO__Y6 $T=502265 106895 0 0 $X=502265 $Y=106895
X659 11 MASCO__Y6 $T=502265 111895 0 0 $X=502265 $Y=111895
X660 11 MASCO__Y6 $T=502265 116895 0 0 $X=502265 $Y=116895
X661 11 MASCO__Y6 $T=502265 121895 0 0 $X=502265 $Y=121895
X662 11 MASCO__Y6 $T=502265 126895 0 0 $X=502265 $Y=126895
X663 11 MASCO__Y6 $T=502265 131895 0 0 $X=502265 $Y=131895
X664 11 MASCO__Y6 $T=502265 136895 0 0 $X=502265 $Y=136895
X665 11 MASCO__Y6 $T=502265 141895 0 0 $X=502265 $Y=141895
X666 11 MASCO__Y6 $T=520265 51895 0 0 $X=520265 $Y=51895
X667 11 MASCO__Y6 $T=520265 56895 0 0 $X=520265 $Y=56895
X668 11 MASCO__Y6 $T=520265 61895 0 0 $X=520265 $Y=61895
X669 11 MASCO__Y6 $T=520265 66895 0 0 $X=520265 $Y=66895
X670 11 MASCO__Y6 $T=520265 71895 0 0 $X=520265 $Y=71895
X671 11 MASCO__Y6 $T=520265 76895 0 0 $X=520265 $Y=76895
X672 11 MASCO__Y6 $T=520265 81895 0 0 $X=520265 $Y=81895
X673 11 MASCO__Y6 $T=520265 86895 0 0 $X=520265 $Y=86895
X674 11 MASCO__Y6 $T=520265 91895 0 0 $X=520265 $Y=91895
X675 11 MASCO__Y6 $T=520265 96895 0 0 $X=520265 $Y=96895
X676 11 MASCO__Y6 $T=520265 101895 0 0 $X=520265 $Y=101895
X677 11 MASCO__Y6 $T=520265 106895 0 0 $X=520265 $Y=106895
X678 11 MASCO__Y6 $T=520265 111895 0 0 $X=520265 $Y=111895
X679 11 MASCO__Y6 $T=520265 116895 0 0 $X=520265 $Y=116895
X680 11 MASCO__Y6 $T=520265 121895 0 0 $X=520265 $Y=121895
X681 11 MASCO__Y6 $T=520265 126895 0 0 $X=520265 $Y=126895
X682 11 MASCO__Y6 $T=520265 131895 0 0 $X=520265 $Y=131895
X683 11 MASCO__Y6 $T=520265 136895 0 0 $X=520265 $Y=136895
X684 11 MASCO__Y6 $T=520265 141895 0 0 $X=520265 $Y=141895
X685 11 MASCO__Y6 $T=538265 51895 0 0 $X=538265 $Y=51895
X686 11 MASCO__Y6 $T=538265 56895 0 0 $X=538265 $Y=56895
X687 11 MASCO__Y6 $T=538265 61895 0 0 $X=538265 $Y=61895
X688 11 MASCO__Y6 $T=538265 66895 0 0 $X=538265 $Y=66895
X689 11 MASCO__Y6 $T=538265 71895 0 0 $X=538265 $Y=71895
X690 11 MASCO__Y6 $T=538265 76895 0 0 $X=538265 $Y=76895
X691 11 MASCO__Y6 $T=538265 81895 0 0 $X=538265 $Y=81895
X692 11 MASCO__Y6 $T=538265 86895 0 0 $X=538265 $Y=86895
X693 11 MASCO__Y6 $T=538265 91895 0 0 $X=538265 $Y=91895
X694 11 MASCO__Y6 $T=538265 96895 0 0 $X=538265 $Y=96895
X695 11 MASCO__Y6 $T=538265 101895 0 0 $X=538265 $Y=101895
X696 11 MASCO__Y6 $T=538265 106895 0 0 $X=538265 $Y=106895
X697 11 MASCO__Y6 $T=538265 111895 0 0 $X=538265 $Y=111895
X698 11 MASCO__Y6 $T=538265 116895 0 0 $X=538265 $Y=116895
X699 11 MASCO__Y6 $T=538265 121895 0 0 $X=538265 $Y=121895
X700 11 MASCO__Y6 $T=538265 126895 0 0 $X=538265 $Y=126895
X701 11 MASCO__Y6 $T=538265 131895 0 0 $X=538265 $Y=131895
X702 11 MASCO__Y6 $T=538265 136895 0 0 $X=538265 $Y=136895
X703 11 MASCO__Y6 $T=538265 141895 0 0 $X=538265 $Y=141895
X704 7 MASCO__Y7 $T=377695 52895 0 0 $X=377695 $Y=52895
X705 7 MASCO__Y7 $T=377695 76895 0 0 $X=377695 $Y=76895
X706 7 MASCO__Y7 $T=377695 100895 0 0 $X=377695 $Y=100895
X707 7 MASCO__Y7 $T=391695 52895 0 0 $X=391695 $Y=52895
X708 7 MASCO__Y7 $T=391695 76895 0 0 $X=391695 $Y=76895
X709 7 MASCO__Y7 $T=391695 100895 0 0 $X=391695 $Y=100895
X710 7 MASCO__Y7 $T=405695 52895 0 0 $X=405695 $Y=52895
X711 7 MASCO__Y7 $T=405695 76895 0 0 $X=405695 $Y=76895
X712 7 MASCO__Y7 $T=405695 100895 0 0 $X=405695 $Y=100895
X713 7 MASCO__Y7 $T=419695 52895 0 0 $X=419695 $Y=52895
X714 7 MASCO__Y7 $T=419695 76895 0 0 $X=419695 $Y=76895
X715 7 MASCO__Y7 $T=419695 100895 0 0 $X=419695 $Y=100895
X716 11 MASCO__Y7 $T=501265 52895 0 0 $X=501265 $Y=52895
X717 11 MASCO__Y7 $T=501265 76895 0 0 $X=501265 $Y=76895
X718 11 MASCO__Y7 $T=501265 100895 0 0 $X=501265 $Y=100895
X719 11 MASCO__Y7 $T=515265 52895 0 0 $X=515265 $Y=52895
X720 11 MASCO__Y7 $T=515265 76895 0 0 $X=515265 $Y=76895
X721 11 MASCO__Y7 $T=515265 100895 0 0 $X=515265 $Y=100895
X722 11 MASCO__Y7 $T=529265 52895 0 0 $X=529265 $Y=52895
X723 11 MASCO__Y7 $T=529265 76895 0 0 $X=529265 $Y=76895
X724 11 MASCO__Y7 $T=529265 100895 0 0 $X=529265 $Y=100895
X725 11 MASCO__Y7 $T=543265 52895 0 0 $X=543265 $Y=52895
X726 11 MASCO__Y7 $T=543265 76895 0 0 $X=543265 $Y=76895
X727 11 MASCO__Y7 $T=543265 100895 0 0 $X=543265 $Y=100895
X728 7 MASCO__Y8 $T=377695 124895 0 0 $X=377695 $Y=124895
X729 7 MASCO__Y8 $T=391695 124895 0 0 $X=391695 $Y=124895
X730 7 MASCO__Y8 $T=405695 124895 0 0 $X=405695 $Y=124895
X731 7 MASCO__Y8 $T=419695 124895 0 0 $X=419695 $Y=124895
X732 11 MASCO__Y8 $T=501265 124895 0 0 $X=501265 $Y=124895
X733 11 MASCO__Y8 $T=515265 124895 0 0 $X=515265 $Y=124895
X734 11 MASCO__Y8 $T=529265 124895 0 0 $X=529265 $Y=124895
X735 11 MASCO__Y8 $T=543265 124895 0 0 $X=543265 $Y=124895
X736 7 MASCO__Y9 $T=377695 50835 0 0 $X=377695 $Y=50835
X737 7 MASCO__Y9 $T=377695 146895 0 0 $X=377695 $Y=146895
X738 7 MASCO__Y9 $T=388695 50835 0 0 $X=388695 $Y=50835
X739 7 MASCO__Y9 $T=388695 146895 0 0 $X=388695 $Y=146895
X740 7 MASCO__Y9 $T=399695 50835 0 0 $X=399695 $Y=50835
X741 7 MASCO__Y9 $T=399695 146895 0 0 $X=399695 $Y=146895
X742 7 MASCO__Y9 $T=410695 50835 0 0 $X=410695 $Y=50835
X743 7 MASCO__Y9 $T=410695 146895 0 0 $X=410695 $Y=146895
X744 7 MASCO__Y9 $T=421695 50835 0 0 $X=421695 $Y=50835
X745 7 MASCO__Y9 $T=421695 146895 0 0 $X=421695 $Y=146895
X746 11 MASCO__Y9 $T=501265 50835 0 0 $X=501265 $Y=50835
X747 11 MASCO__Y9 $T=501265 146895 0 0 $X=501265 $Y=146895
X748 11 MASCO__Y9 $T=512265 50835 0 0 $X=512265 $Y=50835
X749 11 MASCO__Y9 $T=512265 146895 0 0 $X=512265 $Y=146895
X750 11 MASCO__Y9 $T=523265 50835 0 0 $X=523265 $Y=50835
X751 11 MASCO__Y9 $T=523265 146895 0 0 $X=523265 $Y=146895
X752 11 MASCO__Y9 $T=534265 50835 0 0 $X=534265 $Y=50835
X753 11 MASCO__Y9 $T=534265 146895 0 0 $X=534265 $Y=146895
X754 11 MASCO__Y9 $T=545265 50835 0 0 $X=545265 $Y=50835
X755 11 MASCO__Y9 $T=545265 146895 0 0 $X=545265 $Y=146895
X756 2 1 1 MOSVC3 w=2e-05 l=3e-05 $X=16180 $Y=110530 $dt=4
X757 2 1 1 MOSVC3 w=2e-05 l=3e-05 $X=16180 $Y=132530 $dt=4
X758 2 1 1 MOSVC3 w=2e-05 l=3e-05 $X=48780 $Y=110530 $dt=4
X759 2 1 1 MOSVC3 w=2e-05 l=3e-05 $X=48780 $Y=132530 $dt=4
D4 1 2 p_dnw AREA=3.57048e-11 PJ=3.588e-05 perimeter=3.588e-05 $X=11740 $Y=84695 $dt=6
D5 1 2 p_dnw AREA=1.90124e-10 PJ=7.516e-05 perimeter=7.516e-05 $X=59815 $Y=81480 $dt=6
D6 1 2 p_dnw AREA=1.58288e-09 PJ=0.00049318 perimeter=0.00049318 $X=99710 $Y=59910 $dt=6
D7 1 2 p_dnw AREA=3.09086e-09 PJ=0.00032604 perimeter=0.00032604 $X=101390 $Y=114415 $dt=6
D8 1 17 p_dnw AREA=1.82058e-10 PJ=5.826e-05 perimeter=5.826e-05 $X=105905 $Y=15300 $dt=6
D9 1 18 p_dnw AREA=1.82058e-10 PJ=5.826e-05 perimeter=5.826e-05 $X=105905 $Y=44920 $dt=6
D10 1 18 p_dnw AREA=1.82058e-10 PJ=5.826e-05 perimeter=5.826e-05 $X=160185 $Y=15300 $dt=6
D11 1 17 p_dnw AREA=1.82058e-10 PJ=5.826e-05 perimeter=5.826e-05 $X=160185 $Y=44920 $dt=6
D12 1 2 p_dnw AREA=8.36476e-09 PJ=0.0003905 perimeter=0.0003905 $X=226790 $Y=95600 $dt=6
D13 1 2 p_dnw3 AREA=4.20992e-11 PJ=0 perimeter=0 $X=12880 $Y=85835 $dt=9
D14 1 1 p_dnw3 AREA=5.9176e-11 PJ=0.00010492 perimeter=0.00010492 $X=15380 $Y=110100 $dt=9
D15 1 1 p_dnw3 AREA=5.9176e-11 PJ=0.00010492 perimeter=0.00010492 $X=15380 $Y=132100 $dt=9
D16 1 1 p_dnw3 AREA=5.9176e-11 PJ=0.00010492 perimeter=0.00010492 $X=47980 $Y=110100 $dt=9
D17 1 1 p_dnw3 AREA=5.9176e-11 PJ=0.00010492 perimeter=0.00010492 $X=47980 $Y=132100 $dt=9
D18 1 2 p_dnw3 AREA=1.56539e-10 PJ=0 perimeter=0 $X=61455 $Y=83900 $dt=9
D19 1 17 p_dnw3 AREA=5.86064e-10 PJ=7.406e-05 perimeter=7.406e-05 $X=105905 $Y=18860 $dt=9
D20 1 18 p_dnw3 AREA=5.86064e-10 PJ=7.406e-05 perimeter=7.406e-05 $X=105905 $Y=33460 $dt=9
D21 1 2 p_dnw3 AREA=1.22554e-09 PJ=0 perimeter=0 $X=108190 $Y=68670 $dt=9
D22 1 2 p_dnw3 AREA=1.15225e-09 PJ=0.00012214 perimeter=0.00012214 $X=108190 $Y=82290 $dt=9
D23 1 2 p_dnw3 AREA=1.15028e-09 PJ=0 perimeter=0 $X=112150 $Y=124955 $dt=9
D24 1 2 p_dnw3 AREA=1.15028e-09 PJ=0 perimeter=0 $X=112150 $Y=137935 $dt=9
D25 1 18 p_dnw3 AREA=5.86064e-10 PJ=7.406e-05 perimeter=7.406e-05 $X=160185 $Y=18860 $dt=9
D26 1 17 p_dnw3 AREA=5.86064e-10 PJ=7.406e-05 perimeter=7.406e-05 $X=160185 $Y=33460 $dt=9
C27 20 27 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=231620 $Y=128940 $dt=12
C28 20 27 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=263220 $Y=97740 $dt=12
C29 20 27 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=263220 $Y=128940 $dt=12
C30 20 27 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=294820 $Y=97740 $dt=12
C31 20 27 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=294820 $Y=128940 $dt=12
C32 20 27 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=326420 $Y=97740 $dt=12
C33 20 27 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=326420 $Y=128940 $dt=12
.ends current_source_gm_10_en_r

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: mosvc3_CDNS_7246548160521                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt mosvc3_CDNS_7246548160521 1 2
** N=2 EP=2 FDC=2
X0 2 1 1 MOSVC3 w=2.5e-05 l=2e-05 $X=0 $Y=0 $dt=4
D1 1 1 p_dnw3 AREA=5.8576e-11 PJ=9.492e-05 perimeter=9.492e-05 $X=-800 $Y=-430 $dt=9
.ends mosvc3_CDNS_7246548160521

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: mosvc3_CDNS_7246548160522                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt mosvc3_CDNS_7246548160522 1 2
** N=2 EP=2 FDC=2
X0 2 1 1 MOSVC3 w=2e-05 l=2e-05 $X=0 $Y=0 $dt=4
D1 1 1 p_dnw3 AREA=5.0576e-11 PJ=8.492e-05 perimeter=8.492e-05 $X=-800 $Y=-430 $dt=9
.ends mosvc3_CDNS_7246548160522

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160558                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160558 1 2
** N=2 EP=2 FDC=0
.ends VIA1_C_CDNS_7246548160558

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160559                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160559 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246548160559

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160560                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160560 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246548160560

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160561                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160561 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246548160561

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160562                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160562 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246548160562

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246548160563                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246548160563 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246548160563

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160564                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160564 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246548160564

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246548160565                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246548160565 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246548160565

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160567                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160567 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246548160567

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246548160568                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246548160568 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246548160568

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160569                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160569 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246548160569

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_7246548160570                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_7246548160570 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_7246548160570

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246548160571                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246548160571 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246548160571

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160573                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160573 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246548160573

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246548160574                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246548160574 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246548160574

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160575                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160575 1 2
** N=2 EP=2 FDC=0
.ends VIA1_C_CDNS_7246548160575

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246548160576                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246548160576 1 2
** N=2 EP=2 FDC=0
.ends VIA2_C_CDNS_7246548160576

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160577                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160577 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246548160577

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246548160580                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246548160580 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246548160580

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246548160581                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246548160581 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246548160581

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_7246548160584                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_7246548160584 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_7246548160584

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_7246548160586                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_7246548160586 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_7246548160586

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246548160588                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246548160588 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246548160588

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160523                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160523 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
M0 3 2 1 1 pe3 L=1e-05 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
.ends pe3_CDNS_7246548160523

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160524                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160524 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=2
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=2
.ends pe3_CDNS_7246548160524

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160525                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160525 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=4
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=2
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=2
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=2
.ends pe3_CDNS_7246548160525

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160526                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160526 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=8
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=2
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=2
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=2
M4 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=6160 $Y=0 $dt=2
M5 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7700 $Y=0 $dt=2
M6 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=9240 $Y=0 $dt=2
M7 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=10780 $Y=0 $dt=2
.ends pe3_CDNS_7246548160526

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160527                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160527 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=16
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=2
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=2
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=2
M4 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=6160 $Y=0 $dt=2
M5 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7700 $Y=0 $dt=2
M6 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=9240 $Y=0 $dt=2
M7 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10780 $Y=0 $dt=2
M8 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12320 $Y=0 $dt=2
M9 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=13860 $Y=0 $dt=2
M10 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=15400 $Y=0 $dt=2
M11 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=16940 $Y=0 $dt=2
M12 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=18480 $Y=0 $dt=2
M13 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=20020 $Y=0 $dt=2
M14 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=21560 $Y=0 $dt=2
M15 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=23100 $Y=0 $dt=2
.ends pe3_CDNS_7246548160527

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160528                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160528 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=32
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=2
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=2
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=2
M4 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=6160 $Y=0 $dt=2
M5 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7700 $Y=0 $dt=2
M6 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=9240 $Y=0 $dt=2
M7 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10780 $Y=0 $dt=2
M8 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12320 $Y=0 $dt=2
M9 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=13860 $Y=0 $dt=2
M10 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=15400 $Y=0 $dt=2
M11 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=16940 $Y=0 $dt=2
M12 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=18480 $Y=0 $dt=2
M13 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=20020 $Y=0 $dt=2
M14 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=21560 $Y=0 $dt=2
M15 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=23100 $Y=0 $dt=2
M16 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=24640 $Y=0 $dt=2
M17 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=26180 $Y=0 $dt=2
M18 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=27720 $Y=0 $dt=2
M19 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=29260 $Y=0 $dt=2
M20 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=30800 $Y=0 $dt=2
M21 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=32340 $Y=0 $dt=2
M22 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=33880 $Y=0 $dt=2
M23 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=35420 $Y=0 $dt=2
M24 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=36960 $Y=0 $dt=2
M25 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=38500 $Y=0 $dt=2
M26 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=40040 $Y=0 $dt=2
M27 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=41580 $Y=0 $dt=2
M28 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=43120 $Y=0 $dt=2
M29 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=44660 $Y=0 $dt=2
M30 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=46200 $Y=0 $dt=2
M31 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=47740 $Y=0 $dt=2
.ends pe3_CDNS_7246548160528

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7246548160529                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7246548160529 1 2
** N=2 EP=2 FDC=1
R0 2 1 L=0.00021702 W=4e-06 $[rpp1k1_3] $SUB=2 $X=-4220 $Y=0 $dt=10
.ends rpp1k1_3_CDNS_7246548160529

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160530                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160530 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=10
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=2
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=2
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=2
M4 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=6160 $Y=0 $dt=2
M5 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7700 $Y=0 $dt=2
M6 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=9240 $Y=0 $dt=2
M7 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10780 $Y=0 $dt=2
M8 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12320 $Y=0 $dt=2
M9 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=13860 $Y=0 $dt=2
.ends pe3_CDNS_7246548160530

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7246548160531                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7246548160531 1 2
** N=2 EP=2 FDC=1
R0 2 1 L=0.0008227 W=4e-06 $[rpp1k1_3] $SUB=2 $X=-4220 $Y=0 $dt=10
.ends rpp1k1_3_CDNS_7246548160531

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160532                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160532 1 2 3
*.DEVICECLIMB
** N=3 EP=3 FDC=1
M0 2 2 1 1 pe3 L=2e-05 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
.ends pe3_CDNS_7246548160532

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160533                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160533 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
M0 3 2 1 1 pe3 L=3e-07 W=6e-06 AD=2.88e-12 AS=2.88e-12 PD=1.296e-05 PS=1.296e-05 $X=0 $Y=0 $dt=2
.ends pe3_CDNS_7246548160533

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160534                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160534 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=2
M0 3 2 1 4 pe3 L=3.5e-07 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
M1 1 2 3 4 pe3 L=3.5e-07 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=890 $Y=0 $dt=2
.ends pe3_CDNS_7246548160534

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7246548160535                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7246548160535 1 2 3 4
** N=4 EP=4 FDC=8
M0 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=2540 $Y=0 $dt=1
M2 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=5080 $Y=0 $dt=1
M3 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7620 $Y=0 $dt=1
M4 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10160 $Y=0 $dt=1
M5 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12700 $Y=0 $dt=1
M6 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=15240 $Y=0 $dt=1
M7 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=17780 $Y=0 $dt=1
.ends ne3_CDNS_7246548160535

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3i_6_CDNS_7246548160536                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3i_6_CDNS_7246548160536 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=1
X0 1 2 3 1 4 5 NE3I_6 w=1e-05 l=2e-06 as=4.8e-12 ad=4.8e-12 ps=2.096e-05 pd=2.096e-05 $X=0 $Y=0 $dt=3
.ends ne3i_6_CDNS_7246548160536

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7246548160537                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7246548160537 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=2e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends ne3_CDNS_7246548160537

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246548160538                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246548160538 1 2
*.DEVICECLIMB
** N=2 EP=2 FDC=1
M0 1 1 1 1 pe3 L=1e-05 W=2e-06 AD=9.6e-13 AS=9.6e-13 PD=4.96e-06 PS=4.96e-06 $X=0 $Y=0 $dt=2
.ends pe3_CDNS_7246548160538

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7246548160539                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7246548160539 1 2 3
** N=3 EP=3 FDC=4
M0 3 2 1 1 ne3 L=3.5e-07 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 1 ne3 L=3.5e-07 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=890 $Y=0 $dt=1
M2 3 2 1 1 ne3 L=3.5e-07 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1780 $Y=0 $dt=1
M3 1 2 3 1 ne3 L=3.5e-07 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=2670 $Y=0 $dt=1
.ends ne3_CDNS_7246548160539

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A15                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A15 1 2 3 4 5 6 7 8
*.DEVICECLIMB
** N=8 EP=8 FDC=4
X0 3 2 1 8 pe3_CDNS_7246548160523 $T=1510 11030 1 0 $X=0 $Y=0
X1 3 5 4 8 pe3_CDNS_7246548160523 $T=12750 11030 1 0 $X=11240 $Y=0
X2 3 5 6 8 pe3_CDNS_7246548160523 $T=23990 11030 1 0 $X=22480 $Y=0
X3 3 5 7 8 pe3_CDNS_7246548160523 $T=35230 11030 1 0 $X=33720 $Y=0
.ends MASCO__A15

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: dac6b_amp_n2                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt dac6b_amp_n2 1 2 3 4 5 6 7 8 9 10
+ 11 12
** N=31 EP=12 FDC=372
X0 13 VIA1_C_CDNS_724654816055 $T=7445 56365 0 0 $X=7045 $Y=55655
X1 3 VIA1_C_CDNS_724654816055 $T=9985 58145 0 0 $X=9585 $Y=57435
X2 13 VIA1_C_CDNS_724654816055 $T=12525 56365 0 0 $X=12125 $Y=55655
X3 3 VIA1_C_CDNS_724654816055 $T=15065 58145 0 0 $X=14665 $Y=57435
X4 13 VIA1_C_CDNS_724654816055 $T=17605 56365 0 0 $X=17205 $Y=55655
X5 3 VIA1_C_CDNS_724654816055 $T=20145 58145 0 0 $X=19745 $Y=57435
X6 13 VIA1_C_CDNS_724654816055 $T=22685 56365 0 0 $X=22285 $Y=55655
X7 3 VIA1_C_CDNS_724654816055 $T=25225 58145 0 0 $X=24825 $Y=57435
X8 13 VIA1_C_CDNS_724654816055 $T=27765 56365 0 0 $X=27365 $Y=55655
X9 14 VIA1_C_CDNS_724654816055 $T=34200 58145 0 0 $X=33800 $Y=57435
X10 15 VIA1_C_CDNS_724654816055 $T=36740 56365 0 0 $X=36340 $Y=55655
X11 14 VIA1_C_CDNS_724654816055 $T=39280 58145 0 0 $X=38880 $Y=57435
X12 15 VIA1_C_CDNS_724654816055 $T=41820 56365 0 0 $X=41420 $Y=55655
X13 14 VIA1_C_CDNS_724654816055 $T=44360 58145 0 0 $X=43960 $Y=57435
X14 15 VIA1_C_CDNS_724654816055 $T=46900 56365 0 0 $X=46500 $Y=55655
X15 14 VIA1_C_CDNS_724654816055 $T=49440 58145 0 0 $X=49040 $Y=57435
X16 15 VIA1_C_CDNS_724654816055 $T=51980 56365 0 0 $X=51580 $Y=55655
X17 14 VIA1_C_CDNS_724654816055 $T=54520 58145 0 0 $X=54120 $Y=57435
X18 2 VIA1_C_CDNS_724654816055 $T=56070 146660 0 0 $X=55670 $Y=145950
X19 2 VIA1_C_CDNS_724654816055 $T=56070 173480 0 0 $X=55670 $Y=172770
X20 2 VIA1_C_CDNS_724654816055 $T=66380 146660 0 0 $X=65980 $Y=145950
X21 2 VIA1_C_CDNS_724654816055 $T=66380 173480 0 0 $X=65980 $Y=172770
X22 2 VIA1_C_CDNS_724654816055 $T=67540 146660 0 0 $X=67140 $Y=145950
X23 2 VIA1_C_CDNS_724654816055 $T=67540 173480 0 0 $X=67140 $Y=172770
X24 16 VIA1_C_CDNS_724654816055 $T=77620 144880 0 0 $X=77220 $Y=144170
X25 17 VIA1_C_CDNS_724654816055 $T=77620 175260 0 0 $X=77220 $Y=174550
X26 17 VIA1_C_CDNS_724654816055 $T=88860 143100 0 0 $X=88460 $Y=142390
X27 16 VIA1_C_CDNS_724654816055 $T=88860 177040 0 0 $X=88460 $Y=176330
X28 16 VIA1_C_CDNS_724654816055 $T=100100 144880 0 0 $X=99700 $Y=144170
X29 17 VIA1_C_CDNS_724654816055 $T=100100 175260 0 0 $X=99700 $Y=174550
X30 17 VIA1_C_CDNS_724654816055 $T=111340 143100 0 0 $X=110940 $Y=142390
X31 16 VIA1_C_CDNS_724654816055 $T=111340 177040 0 0 $X=110940 $Y=176330
X32 16 VIA1_C_CDNS_724654816055 $T=122580 144880 0 0 $X=122180 $Y=144170
X33 17 VIA1_C_CDNS_724654816055 $T=122580 175260 0 0 $X=122180 $Y=174550
X34 17 VIA1_C_CDNS_724654816055 $T=133820 143100 0 0 $X=133420 $Y=142390
X35 16 VIA1_C_CDNS_724654816055 $T=133820 177040 0 0 $X=133420 $Y=176330
X36 16 VIA1_C_CDNS_724654816055 $T=145060 144880 0 0 $X=144660 $Y=144170
X37 17 VIA1_C_CDNS_724654816055 $T=145060 175260 0 0 $X=144660 $Y=174550
X38 18 VIA1_C_CDNS_724654816055 $T=154405 72995 0 0 $X=154005 $Y=72285
X39 19 VIA1_C_CDNS_724654816055 $T=154405 94475 0 0 $X=154005 $Y=93765
X40 20 VIA1_C_CDNS_724654816055 $T=154405 115425 0 0 $X=154005 $Y=114715
X41 17 VIA1_C_CDNS_724654816055 $T=156300 143100 0 0 $X=155900 $Y=142390
X42 16 VIA1_C_CDNS_724654816055 $T=156300 177040 0 0 $X=155900 $Y=176330
X43 2 VIA1_C_CDNS_724654816055 $T=167770 146660 0 0 $X=167370 $Y=145950
X44 2 VIA1_C_CDNS_724654816055 $T=167770 173480 0 0 $X=167370 $Y=172770
X45 1 VIA1_C_CDNS_724654816055 $T=174945 74775 0 0 $X=174545 $Y=74065
X46 18 VIA1_C_CDNS_724654816055 $T=174945 96255 0 0 $X=174545 $Y=95545
X47 19 VIA1_C_CDNS_724654816055 $T=174945 117205 0 0 $X=174545 $Y=116495
X48 21 VIA1_C_CDNS_724654816056 $T=61935 55475 0 0 $X=61795 $Y=54505
X49 22 VIA1_C_CDNS_724654816056 $T=64475 57755 0 0 $X=64335 $Y=56785
X50 21 VIA1_C_CDNS_724654816056 $T=67015 55475 0 0 $X=66875 $Y=54505
X51 22 VIA1_C_CDNS_724654816056 $T=69555 57755 0 0 $X=69415 $Y=56785
X52 21 VIA1_C_CDNS_724654816056 $T=72095 55475 0 0 $X=71955 $Y=54505
X53 22 VIA1_C_CDNS_724654816056 $T=74635 57755 0 0 $X=74495 $Y=56785
X54 21 VIA1_C_CDNS_724654816056 $T=77175 55475 0 0 $X=77035 $Y=54505
X55 22 VIA1_C_CDNS_724654816056 $T=79715 57755 0 0 $X=79575 $Y=56785
X56 21 VIA1_C_CDNS_724654816056 $T=82255 55475 0 0 $X=82115 $Y=54505
X57 3 VIA1_C_CDNS_724654816057 $T=8715 70535 0 0 $X=8315 $Y=70345
X58 3 VIA1_C_CDNS_724654816057 $T=11255 70535 0 0 $X=10855 $Y=70345
X59 3 VIA1_C_CDNS_724654816057 $T=13795 70535 0 0 $X=13395 $Y=70345
X60 13 VIA1_C_CDNS_724654816057 $T=15770 27420 0 0 $X=15370 $Y=27230
X61 3 VIA1_C_CDNS_724654816057 $T=16335 70535 0 0 $X=15935 $Y=70345
X62 3 VIA1_C_CDNS_724654816057 $T=18875 70535 0 0 $X=18475 $Y=70345
X63 13 VIA1_C_CDNS_724654816057 $T=19010 27420 0 0 $X=18610 $Y=27230
X64 15 VIA1_C_CDNS_724654816057 $T=20710 160140 0 0 $X=20310 $Y=159950
X65 3 VIA1_C_CDNS_724654816057 $T=21415 70535 0 0 $X=21015 $Y=70345
X66 13 VIA1_C_CDNS_724654816057 $T=22250 27420 0 0 $X=21850 $Y=27230
X67 3 VIA1_C_CDNS_724654816057 $T=23955 70535 0 0 $X=23555 $Y=70345
X68 13 VIA1_C_CDNS_724654816057 $T=25490 27420 0 0 $X=25090 $Y=27230
X69 3 VIA1_C_CDNS_724654816057 $T=26495 70535 0 0 $X=26095 $Y=70345
X70 13 VIA1_C_CDNS_724654816057 $T=28730 27420 0 0 $X=28330 $Y=27230
X71 15 VIA1_C_CDNS_724654816057 $T=31950 160140 0 0 $X=31550 $Y=159950
X72 13 VIA1_C_CDNS_724654816057 $T=31970 27420 0 0 $X=31570 $Y=27230
X73 13 VIA1_C_CDNS_724654816057 $T=35210 27420 0 0 $X=34810 $Y=27230
X74 3 VIA1_C_CDNS_724654816057 $T=35470 70535 0 0 $X=35070 $Y=70345
X75 3 VIA1_C_CDNS_724654816057 $T=38010 70535 0 0 $X=37610 $Y=70345
X76 13 VIA1_C_CDNS_724654816057 $T=38450 27420 0 0 $X=38050 $Y=27230
X77 3 VIA1_C_CDNS_724654816057 $T=40550 70535 0 0 $X=40150 $Y=70345
X78 13 VIA1_C_CDNS_724654816057 $T=41690 27420 0 0 $X=41290 $Y=27230
X79 3 VIA1_C_CDNS_724654816057 $T=43090 70535 0 0 $X=42690 $Y=70345
X80 13 VIA1_C_CDNS_724654816057 $T=44930 27420 0 0 $X=44530 $Y=27230
X81 3 VIA1_C_CDNS_724654816057 $T=45630 70535 0 0 $X=45230 $Y=70345
X82 13 VIA1_C_CDNS_724654816057 $T=48170 27420 0 0 $X=47770 $Y=27230
X83 3 VIA1_C_CDNS_724654816057 $T=48170 70535 0 0 $X=47770 $Y=70345
X84 3 VIA1_C_CDNS_724654816057 $T=50710 70535 0 0 $X=50310 $Y=70345
X85 13 VIA1_C_CDNS_724654816057 $T=51410 27420 0 0 $X=51010 $Y=27230
X86 3 VIA1_C_CDNS_724654816057 $T=53250 70535 0 0 $X=52850 $Y=70345
X87 3 VIA1_C_CDNS_724654816057 $T=63205 70535 0 0 $X=62805 $Y=70345
X88 3 VIA1_C_CDNS_724654816057 $T=65745 70535 0 0 $X=65345 $Y=70345
X89 3 VIA1_C_CDNS_724654816057 $T=68285 70535 0 0 $X=67885 $Y=70345
X90 3 VIA1_C_CDNS_724654816057 $T=70825 70535 0 0 $X=70425 $Y=70345
X91 16 VIA1_C_CDNS_724654816057 $T=72580 160140 0 0 $X=72180 $Y=159950
X92 3 VIA1_C_CDNS_724654816057 $T=73365 70535 0 0 $X=72965 $Y=70345
X93 3 VIA1_C_CDNS_724654816057 $T=75905 70535 0 0 $X=75505 $Y=70345
X94 3 VIA1_C_CDNS_724654816057 $T=78445 70535 0 0 $X=78045 $Y=70345
X95 3 VIA1_C_CDNS_724654816057 $T=80985 70535 0 0 $X=80585 $Y=70345
X96 16 VIA1_C_CDNS_724654816057 $T=83820 160140 0 0 $X=83420 $Y=159950
X97 16 VIA1_C_CDNS_724654816057 $T=95060 160140 0 0 $X=94660 $Y=159950
X98 16 VIA1_C_CDNS_724654816057 $T=106300 160140 0 0 $X=105900 $Y=159950
X99 16 VIA1_C_CDNS_724654816057 $T=117540 160140 0 0 $X=117140 $Y=159950
X100 16 VIA1_C_CDNS_724654816057 $T=128780 160140 0 0 $X=128380 $Y=159950
X101 16 VIA1_C_CDNS_724654816057 $T=140020 160140 0 0 $X=139620 $Y=159950
X102 16 VIA1_C_CDNS_724654816057 $T=151260 160140 0 0 $X=150860 $Y=159950
X103 19 VIA1_C_CDNS_724654816057 $T=224435 24760 0 0 $X=224035 $Y=24570
X104 19 VIA1_C_CDNS_724654816057 $T=225975 24760 0 0 $X=225575 $Y=24570
X105 19 VIA1_C_CDNS_724654816057 $T=227515 24760 0 0 $X=227115 $Y=24570
X106 19 VIA1_C_CDNS_724654816057 $T=229055 24760 0 0 $X=228655 $Y=24570
X107 19 VIA1_C_CDNS_724654816057 $T=230595 24760 0 0 $X=230195 $Y=24570
X108 19 VIA1_C_CDNS_724654816057 $T=232135 24760 0 0 $X=231735 $Y=24570
X109 19 VIA1_C_CDNS_724654816057 $T=233675 24760 0 0 $X=233275 $Y=24570
X110 19 VIA1_C_CDNS_724654816057 $T=235215 24760 0 0 $X=234815 $Y=24570
X111 19 VIA1_C_CDNS_724654816057 $T=236755 24760 0 0 $X=236355 $Y=24570
X112 19 VIA1_C_CDNS_724654816057 $T=238295 24760 0 0 $X=237895 $Y=24570
X113 19 VIA1_C_CDNS_724654816057 $T=247255 24760 0 0 $X=246855 $Y=24570
X114 19 VIA1_C_CDNS_724654816057 $T=248795 24760 0 0 $X=248395 $Y=24570
X115 19 VIA1_C_CDNS_724654816057 $T=250335 24760 0 0 $X=249935 $Y=24570
X116 19 VIA1_C_CDNS_724654816057 $T=251875 24760 0 0 $X=251475 $Y=24570
X117 19 VIA1_C_CDNS_724654816057 $T=253415 24760 0 0 $X=253015 $Y=24570
X118 19 VIA1_C_CDNS_724654816057 $T=254955 24760 0 0 $X=254555 $Y=24570
X119 19 VIA1_C_CDNS_724654816057 $T=256495 24760 0 0 $X=256095 $Y=24570
X120 19 VIA1_C_CDNS_724654816057 $T=258035 24760 0 0 $X=257635 $Y=24570
X121 19 VIA1_C_CDNS_724654816057 $T=259575 24760 0 0 $X=259175 $Y=24570
X122 19 VIA1_C_CDNS_724654816057 $T=261115 24760 0 0 $X=260715 $Y=24570
X123 19 VIA1_C_CDNS_724654816057 $T=262655 24760 0 0 $X=262255 $Y=24570
X124 19 VIA1_C_CDNS_724654816057 $T=264195 24760 0 0 $X=263795 $Y=24570
X125 19 VIA1_C_CDNS_724654816057 $T=265735 24760 0 0 $X=265335 $Y=24570
X126 19 VIA1_C_CDNS_724654816057 $T=267275 24760 0 0 $X=266875 $Y=24570
X127 19 VIA1_C_CDNS_724654816057 $T=268815 24760 0 0 $X=268415 $Y=24570
X128 19 VIA1_C_CDNS_724654816057 $T=270355 24760 0 0 $X=269955 $Y=24570
X129 19 VIA1_C_CDNS_724654816057 $T=271895 24760 0 0 $X=271495 $Y=24570
X130 19 VIA1_C_CDNS_724654816057 $T=273435 24760 0 0 $X=273035 $Y=24570
X131 19 VIA1_C_CDNS_724654816057 $T=274975 24760 0 0 $X=274575 $Y=24570
X132 19 VIA1_C_CDNS_724654816057 $T=276515 24760 0 0 $X=276115 $Y=24570
X133 19 VIA1_C_CDNS_724654816057 $T=278055 24760 0 0 $X=277655 $Y=24570
X134 19 VIA1_C_CDNS_724654816057 $T=279595 24760 0 0 $X=279195 $Y=24570
X135 19 VIA1_C_CDNS_724654816057 $T=281135 24760 0 0 $X=280735 $Y=24570
X136 19 VIA1_C_CDNS_724654816057 $T=282675 24760 0 0 $X=282275 $Y=24570
X137 19 VIA1_C_CDNS_724654816057 $T=284215 24760 0 0 $X=283815 $Y=24570
X138 19 VIA1_C_CDNS_724654816057 $T=285755 24760 0 0 $X=285355 $Y=24570
X139 19 VIA1_C_CDNS_724654816057 $T=287295 24760 0 0 $X=286895 $Y=24570
X140 19 VIA1_C_CDNS_724654816057 $T=288835 24760 0 0 $X=288435 $Y=24570
X141 19 VIA1_C_CDNS_724654816057 $T=290375 24760 0 0 $X=289975 $Y=24570
X142 19 VIA1_C_CDNS_724654816057 $T=291915 24760 0 0 $X=291515 $Y=24570
X143 19 VIA1_C_CDNS_724654816057 $T=293455 24760 0 0 $X=293055 $Y=24570
X144 19 VIA1_C_CDNS_724654816057 $T=294995 24760 0 0 $X=294595 $Y=24570
X145 19 VIA1_C_CDNS_724654816057 $T=303070 24760 0 0 $X=302670 $Y=24570
X146 19 VIA1_C_CDNS_724654816057 $T=304610 24760 0 0 $X=304210 $Y=24570
X147 19 VIA1_C_CDNS_724654816057 $T=306150 24760 0 0 $X=305750 $Y=24570
X148 19 VIA1_C_CDNS_724654816057 $T=307690 24760 0 0 $X=307290 $Y=24570
X149 19 VIA1_C_CDNS_724654816057 $T=309230 24760 0 0 $X=308830 $Y=24570
X150 19 VIA1_C_CDNS_724654816057 $T=310770 24760 0 0 $X=310370 $Y=24570
X151 19 VIA1_C_CDNS_724654816057 $T=312310 24760 0 0 $X=311910 $Y=24570
X152 19 VIA1_C_CDNS_724654816057 $T=313850 24760 0 0 $X=313450 $Y=24570
X153 19 VIA1_C_CDNS_724654816057 $T=315390 24760 0 0 $X=314990 $Y=24570
X154 19 VIA1_C_CDNS_724654816057 $T=316930 24760 0 0 $X=316530 $Y=24570
X155 19 VIA1_C_CDNS_724654816057 $T=318470 24760 0 0 $X=318070 $Y=24570
X156 19 VIA1_C_CDNS_724654816057 $T=320010 24760 0 0 $X=319610 $Y=24570
X157 19 VIA1_C_CDNS_724654816057 $T=321550 24760 0 0 $X=321150 $Y=24570
X158 19 VIA1_C_CDNS_724654816057 $T=323090 24760 0 0 $X=322690 $Y=24570
X159 19 VIA1_C_CDNS_724654816057 $T=324630 24760 0 0 $X=324230 $Y=24570
X160 19 VIA1_C_CDNS_724654816057 $T=326170 24760 0 0 $X=325770 $Y=24570
X161 19 VIA1_C_CDNS_724654816057 $T=333835 24760 0 0 $X=333435 $Y=24570
X162 19 VIA1_C_CDNS_724654816057 $T=335375 24760 0 0 $X=334975 $Y=24570
X163 19 VIA1_C_CDNS_724654816057 $T=336915 24760 0 0 $X=336515 $Y=24570
X164 19 VIA1_C_CDNS_724654816057 $T=338455 24760 0 0 $X=338055 $Y=24570
X165 19 VIA1_C_CDNS_724654816057 $T=339995 24760 0 0 $X=339595 $Y=24570
X166 19 VIA1_C_CDNS_724654816057 $T=341535 24760 0 0 $X=341135 $Y=24570
X167 19 VIA1_C_CDNS_724654816057 $T=343075 24760 0 0 $X=342675 $Y=24570
X168 19 VIA1_C_CDNS_724654816057 $T=344615 24760 0 0 $X=344215 $Y=24570
X169 19 VIA1_C_CDNS_724654816057 $T=352300 24760 0 0 $X=351900 $Y=24570
X170 19 VIA1_C_CDNS_724654816057 $T=353840 24760 0 0 $X=353440 $Y=24570
X171 19 VIA1_C_CDNS_724654816057 $T=355380 24760 0 0 $X=354980 $Y=24570
X172 19 VIA1_C_CDNS_724654816057 $T=356920 24760 0 0 $X=356520 $Y=24570
X173 19 VIA1_C_CDNS_724654816057 $T=364635 24760 0 0 $X=364235 $Y=24570
X174 19 VIA1_C_CDNS_724654816057 $T=366175 24760 0 0 $X=365775 $Y=24570
X175 19 VIA1_C_CDNS_724654816057 $T=374010 24760 0 0 $X=373610 $Y=24570
X176 13 VIA2_C_CDNS_724654816058 $T=6660 9690 0 0 $X=5690 $Y=9030
X177 13 VIA2_C_CDNS_724654816058 $T=6660 41530 0 0 $X=5690 $Y=40870
X178 16 VIA2_C_CDNS_724654816058 $T=51270 144880 0 0 $X=50300 $Y=144220
X179 16 VIA2_C_CDNS_724654816058 $T=51270 177040 0 0 $X=50300 $Y=176380
X180 14 VIA2_C_CDNS_724654816058 $T=60010 13250 0 0 $X=59040 $Y=12590
X181 14 VIA2_C_CDNS_724654816058 $T=60010 45090 0 0 $X=59040 $Y=44430
X182 21 VIA2_C_CDNS_724654816058 $T=62290 11470 0 0 $X=61320 $Y=10810
X183 21 VIA2_C_CDNS_724654816058 $T=62290 43310 0 0 $X=61320 $Y=42650
X184 17 VIA2_C_CDNS_724654816058 $T=172570 143100 0 0 $X=171600 $Y=142440
X185 17 VIA2_C_CDNS_724654816058 $T=172570 175260 0 0 $X=171600 $Y=174600
X186 13 VIA2_C_CDNS_7246548160510 $T=6660 27420 0 0 $X=5690 $Y=27280
X187 16 VIA2_C_CDNS_7246548160510 $T=51270 160140 0 0 $X=50300 $Y=160000
X188 1 VIA1_C_CDNS_7246548160511 $T=8940 15030 0 0 $X=7970 $Y=14370
X189 1 VIA1_C_CDNS_7246548160511 $T=8940 39750 0 0 $X=7970 $Y=39090
X190 2 VIA1_C_CDNS_7246548160511 $T=12920 146660 0 0 $X=11950 $Y=146000
X191 2 VIA1_C_CDNS_7246548160511 $T=12920 173480 0 0 $X=11950 $Y=172820
X192 2 VIA1_C_CDNS_7246548160511 $T=39740 146660 0 0 $X=38770 $Y=146000
X193 2 VIA1_C_CDNS_7246548160511 $T=39740 173480 0 0 $X=38770 $Y=172820
X194 2 VIA1_C_CDNS_7246548160511 $T=53550 146660 0 0 $X=52580 $Y=146000
X195 2 VIA1_C_CDNS_7246548160511 $T=53550 173480 0 0 $X=52580 $Y=172820
X196 1 VIA1_C_CDNS_7246548160511 $T=57730 15030 0 0 $X=56760 $Y=14370
X197 1 VIA1_C_CDNS_7246548160511 $T=57730 39750 0 0 $X=56760 $Y=39090
X198 2 VIA1_C_CDNS_7246548160511 $T=170290 146660 0 0 $X=169320 $Y=146000
X199 2 VIA1_C_CDNS_7246548160511 $T=170290 173480 0 0 $X=169320 $Y=172820
X200 1 VIA1_C_CDNS_7246548160514 $T=11260 15030 0 0 $X=11120 $Y=14320
X201 1 VIA1_C_CDNS_7246548160514 $T=11260 39750 0 0 $X=11120 $Y=39040
X202 1 VIA1_C_CDNS_7246548160514 $T=13800 15030 0 0 $X=13660 $Y=14320
X203 1 VIA1_C_CDNS_7246548160514 $T=13800 39750 0 0 $X=13660 $Y=39040
X204 1 VIA1_C_CDNS_7246548160514 $T=14500 15030 0 0 $X=14360 $Y=14320
X205 1 VIA1_C_CDNS_7246548160514 $T=14500 39750 0 0 $X=14360 $Y=39040
X206 2 VIA1_C_CDNS_7246548160514 $T=15440 146660 0 0 $X=15300 $Y=145950
X207 2 VIA1_C_CDNS_7246548160514 $T=15440 173480 0 0 $X=15300 $Y=172770
X208 21 VIA1_C_CDNS_7246548160514 $T=17040 11470 0 0 $X=16900 $Y=10760
X209 13 VIA1_C_CDNS_7246548160514 $T=17040 41530 0 0 $X=16900 $Y=40820
X210 1 VIA1_C_CDNS_7246548160514 $T=17740 15030 0 0 $X=17600 $Y=14320
X211 1 VIA1_C_CDNS_7246548160514 $T=17740 39750 0 0 $X=17600 $Y=39040
X212 14 VIA1_C_CDNS_7246548160514 $T=20280 13250 0 0 $X=20140 $Y=12540
X213 21 VIA1_C_CDNS_7246548160514 $T=20280 43310 0 0 $X=20140 $Y=42600
X214 1 VIA1_C_CDNS_7246548160514 $T=20980 15030 0 0 $X=20840 $Y=14320
X215 1 VIA1_C_CDNS_7246548160514 $T=20980 39750 0 0 $X=20840 $Y=39040
X216 13 VIA1_C_CDNS_7246548160514 $T=23520 9690 0 0 $X=23380 $Y=8980
X217 14 VIA1_C_CDNS_7246548160514 $T=23520 45090 0 0 $X=23380 $Y=44380
X218 1 VIA1_C_CDNS_7246548160514 $T=24220 15030 0 0 $X=24080 $Y=14320
X219 1 VIA1_C_CDNS_7246548160514 $T=24220 39750 0 0 $X=24080 $Y=39040
X220 15 VIA1_C_CDNS_7246548160514 $T=25980 144880 0 0 $X=25840 $Y=144170
X221 20 VIA1_C_CDNS_7246548160514 $T=25980 175260 0 0 $X=25840 $Y=174550
X222 2 VIA1_C_CDNS_7246548160514 $T=26680 146660 0 0 $X=26540 $Y=145950
X223 2 VIA1_C_CDNS_7246548160514 $T=26680 173480 0 0 $X=26540 $Y=172770
X224 21 VIA1_C_CDNS_7246548160514 $T=26760 11470 0 0 $X=26620 $Y=10760
X225 13 VIA1_C_CDNS_7246548160514 $T=26760 41530 0 0 $X=26620 $Y=40820
X226 1 VIA1_C_CDNS_7246548160514 $T=27460 15030 0 0 $X=27320 $Y=14320
X227 1 VIA1_C_CDNS_7246548160514 $T=27460 39750 0 0 $X=27320 $Y=39040
X228 14 VIA1_C_CDNS_7246548160514 $T=30000 13250 0 0 $X=29860 $Y=12540
X229 21 VIA1_C_CDNS_7246548160514 $T=30000 43310 0 0 $X=29860 $Y=42600
X230 1 VIA1_C_CDNS_7246548160514 $T=30700 15030 0 0 $X=30560 $Y=14320
X231 1 VIA1_C_CDNS_7246548160514 $T=30700 39750 0 0 $X=30560 $Y=39040
X232 13 VIA1_C_CDNS_7246548160514 $T=33240 9690 0 0 $X=33100 $Y=8980
X233 14 VIA1_C_CDNS_7246548160514 $T=33240 45090 0 0 $X=33100 $Y=44380
X234 1 VIA1_C_CDNS_7246548160514 $T=33940 15030 0 0 $X=33800 $Y=14320
X235 1 VIA1_C_CDNS_7246548160514 $T=33940 39750 0 0 $X=33800 $Y=39040
X236 21 VIA1_C_CDNS_7246548160514 $T=36480 11470 0 0 $X=36340 $Y=10760
X237 13 VIA1_C_CDNS_7246548160514 $T=36480 41530 0 0 $X=36340 $Y=40820
X238 1 VIA1_C_CDNS_7246548160514 $T=37180 15030 0 0 $X=37040 $Y=14320
X239 1 VIA1_C_CDNS_7246548160514 $T=37180 39750 0 0 $X=37040 $Y=39040
X240 20 VIA1_C_CDNS_7246548160514 $T=37220 143100 0 0 $X=37080 $Y=142390
X241 15 VIA1_C_CDNS_7246548160514 $T=37220 177040 0 0 $X=37080 $Y=176330
X242 14 VIA1_C_CDNS_7246548160514 $T=39720 13250 0 0 $X=39580 $Y=12540
X243 21 VIA1_C_CDNS_7246548160514 $T=39720 43310 0 0 $X=39580 $Y=42600
X244 1 VIA1_C_CDNS_7246548160514 $T=40420 15030 0 0 $X=40280 $Y=14320
X245 1 VIA1_C_CDNS_7246548160514 $T=40420 39750 0 0 $X=40280 $Y=39040
X246 13 VIA1_C_CDNS_7246548160514 $T=42960 9690 0 0 $X=42820 $Y=8980
X247 14 VIA1_C_CDNS_7246548160514 $T=42960 45090 0 0 $X=42820 $Y=44380
X248 1 VIA1_C_CDNS_7246548160514 $T=43660 15030 0 0 $X=43520 $Y=14320
X249 1 VIA1_C_CDNS_7246548160514 $T=43660 39750 0 0 $X=43520 $Y=39040
X250 21 VIA1_C_CDNS_7246548160514 $T=46200 11470 0 0 $X=46060 $Y=10760
X251 13 VIA1_C_CDNS_7246548160514 $T=46200 41530 0 0 $X=46060 $Y=40820
X252 1 VIA1_C_CDNS_7246548160514 $T=46900 15030 0 0 $X=46760 $Y=14320
X253 1 VIA1_C_CDNS_7246548160514 $T=46900 39750 0 0 $X=46760 $Y=39040
X254 14 VIA1_C_CDNS_7246548160514 $T=49440 13250 0 0 $X=49300 $Y=12540
X255 21 VIA1_C_CDNS_7246548160514 $T=49440 43310 0 0 $X=49300 $Y=42600
X256 1 VIA1_C_CDNS_7246548160514 $T=50140 15030 0 0 $X=50000 $Y=14320
X257 1 VIA1_C_CDNS_7246548160514 $T=50140 39750 0 0 $X=50000 $Y=39040
X258 13 VIA1_C_CDNS_7246548160514 $T=52680 9690 0 0 $X=52540 $Y=8980
X259 14 VIA1_C_CDNS_7246548160514 $T=52680 45090 0 0 $X=52540 $Y=44380
X260 1 VIA1_C_CDNS_7246548160514 $T=53380 15030 0 0 $X=53240 $Y=14320
X261 1 VIA1_C_CDNS_7246548160514 $T=53380 39750 0 0 $X=53240 $Y=39040
X262 1 VIA1_C_CDNS_7246548160514 $T=55920 15030 0 0 $X=55780 $Y=14320
X263 1 VIA1_C_CDNS_7246548160514 $T=55920 39750 0 0 $X=55780 $Y=39040
X264 4 VIA1_C_CDNS_7246548160519 $T=89720 58980 0 0 $X=88970 $Y=58750
X265 4 VIA1_C_CDNS_7246548160519 $T=89825 61565 0 90 $X=89595 $Y=60815
X266 15 VIA2_C_CDNS_7246548160525 $T=52465 56350 0 0 $X=49895 $Y=55600
X267 5 VIA2_C_CDNS_7246548160535 $T=185295 41010 0 0 $X=184805 $Y=38960
X268 23 VIA1_C_CDNS_7246548160536 $T=75215 41040 0 0 $X=74725 $Y=38990
X269 5 VIA1_C_CDNS_7246548160536 $T=185295 41010 0 0 $X=184805 $Y=38960
X270 2 VIA1_C_CDNS_7246548160539 $T=90930 69330 0 0 $X=88880 $Y=68840
X271 2 VIA1_C_CDNS_7246548160539 $T=90930 73450 0 0 $X=88880 $Y=72960
X272 23 VIA2_C_CDNS_7246548160541 $T=140695 59650 0 0 $X=140465 $Y=57600
X273 4 VIA2_C_CDNS_7246548160543 $T=89070 58460 0 0 $X=88320 $Y=57710
X274 7 VIA2_C_CDNS_7246548160543 $T=307715 6345 0 0 $X=306965 $Y=5595
X275 8 VIA2_C_CDNS_7246548160543 $T=316955 6345 0 0 $X=316205 $Y=5595
X276 9 VIA2_C_CDNS_7246548160543 $T=326225 6345 0 0 $X=325475 $Y=5595
X277 10 VIA2_C_CDNS_7246548160543 $T=335490 6345 0 0 $X=334740 $Y=5595
X278 11 VIA2_C_CDNS_7246548160543 $T=344750 6345 0 0 $X=344000 $Y=5595
X279 12 VIA2_C_CDNS_7246548160543 $T=354005 6345 0 0 $X=353255 $Y=5595
X280 24 19 5 2 1 pe3_CDNS_724654816056 $T=373510 36320 1 0 $X=372000 $Y=25290
X281 1 4 25 ne3_CDNS_7246548160518 $T=91035 56560 0 0 $X=90235 $Y=56160
X282 18 1 VIA1_C_CDNS_7246548160558 $T=166585 72935 0 0 $X=155215 $Y=72795
X283 19 1 VIA1_C_CDNS_7246548160558 $T=166585 94415 0 0 $X=155215 $Y=94275
X284 20 1 VIA1_C_CDNS_7246548160558 $T=166585 115365 0 0 $X=155215 $Y=115225
X285 18 VIA1_C_CDNS_7246548160559 $T=152520 72935 0 0 $X=151290 $Y=72795
X286 19 VIA1_C_CDNS_7246548160559 $T=152520 94415 0 0 $X=151290 $Y=94275
X287 20 VIA1_C_CDNS_7246548160559 $T=152520 115365 0 0 $X=151290 $Y=115225
X288 1 VIA1_C_CDNS_7246548160560 $T=10335 15030 0 0 $X=10195 $Y=14280
X289 1 VIA1_C_CDNS_7246548160560 $T=10335 39750 0 0 $X=10195 $Y=39000
X290 2 VIA1_C_CDNS_7246548160561 $T=214955 116235 0 0 $X=213985 $Y=116095
X291 2 VIA1_C_CDNS_7246548160561 $T=217155 78635 0 0 $X=216185 $Y=78495
X292 2 VIA1_C_CDNS_7246548160561 $T=217155 97435 0 0 $X=216185 $Y=97295
X293 2 VIA1_C_CDNS_7246548160561 $T=217155 116235 0 0 $X=216185 $Y=116095
X294 2 VIA1_C_CDNS_7246548160561 $T=217155 135035 0 0 $X=216185 $Y=134895
X295 2 VIA1_C_CDNS_7246548160561 $T=217155 153835 0 0 $X=216185 $Y=153695
X296 26 VIA1_C_CDNS_7246548160561 $T=226195 114675 0 0 $X=225225 $Y=114535
X297 2 VIA1_C_CDNS_7246548160561 $T=229015 78635 0 0 $X=228045 $Y=78495
X298 2 VIA1_C_CDNS_7246548160561 $T=229015 97435 0 0 $X=228045 $Y=97295
X299 2 VIA1_C_CDNS_7246548160561 $T=229015 116235 0 0 $X=228045 $Y=116095
X300 2 VIA1_C_CDNS_7246548160561 $T=229015 135035 0 0 $X=228045 $Y=134895
X301 2 VIA1_C_CDNS_7246548160561 $T=229015 153835 0 0 $X=228045 $Y=153695
X302 27 VIA1_C_CDNS_7246548160561 $T=237385 113895 0 0 $X=236415 $Y=113755
X303 2 VIA1_C_CDNS_7246548160561 $T=240255 78635 0 0 $X=239285 $Y=78495
X304 2 VIA1_C_CDNS_7246548160561 $T=240255 97435 0 0 $X=239285 $Y=97295
X305 2 VIA1_C_CDNS_7246548160561 $T=240255 116235 0 0 $X=239285 $Y=116095
X306 2 VIA1_C_CDNS_7246548160561 $T=240255 135035 0 0 $X=239285 $Y=134895
X307 2 VIA1_C_CDNS_7246548160561 $T=240255 153835 0 0 $X=239285 $Y=153695
X308 28 VIA1_C_CDNS_7246548160561 $T=248625 113115 0 0 $X=247655 $Y=112975
X309 2 VIA1_C_CDNS_7246548160561 $T=251495 78635 0 0 $X=250525 $Y=78495
X310 2 VIA1_C_CDNS_7246548160561 $T=251495 97435 0 0 $X=250525 $Y=97295
X311 2 VIA1_C_CDNS_7246548160561 $T=251495 116235 0 0 $X=250525 $Y=116095
X312 2 VIA1_C_CDNS_7246548160561 $T=251495 135035 0 0 $X=250525 $Y=134895
X313 2 VIA1_C_CDNS_7246548160561 $T=251495 153835 0 0 $X=250525 $Y=153695
X314 29 VIA1_C_CDNS_7246548160561 $T=259865 111555 0 0 $X=258895 $Y=111415
X315 2 VIA1_C_CDNS_7246548160561 $T=262735 78635 0 0 $X=261765 $Y=78495
X316 2 VIA1_C_CDNS_7246548160561 $T=262735 97435 0 0 $X=261765 $Y=97295
X317 2 VIA1_C_CDNS_7246548160561 $T=262735 116235 0 0 $X=261765 $Y=116095
X318 2 VIA1_C_CDNS_7246548160561 $T=262735 135035 0 0 $X=261765 $Y=134895
X319 2 VIA1_C_CDNS_7246548160561 $T=262735 153835 0 0 $X=261765 $Y=153695
X320 30 VIA1_C_CDNS_7246548160561 $T=271105 115455 0 0 $X=270135 $Y=115315
X321 2 VIA1_C_CDNS_7246548160561 $T=273975 78635 0 0 $X=273005 $Y=78495
X322 2 VIA1_C_CDNS_7246548160561 $T=273975 97435 0 0 $X=273005 $Y=97295
X323 2 VIA1_C_CDNS_7246548160561 $T=273975 116235 0 0 $X=273005 $Y=116095
X324 2 VIA1_C_CDNS_7246548160561 $T=273975 135035 0 0 $X=273005 $Y=134895
X325 2 VIA1_C_CDNS_7246548160561 $T=273975 153835 0 0 $X=273005 $Y=153695
X326 24 VIA1_C_CDNS_7246548160561 $T=282345 109995 0 0 $X=281375 $Y=109855
X327 2 VIA1_C_CDNS_7246548160561 $T=285215 78635 0 0 $X=284245 $Y=78495
X328 2 VIA1_C_CDNS_7246548160561 $T=285215 97435 0 0 $X=284245 $Y=97295
X329 2 VIA1_C_CDNS_7246548160561 $T=285215 116235 0 0 $X=284245 $Y=116095
X330 2 VIA1_C_CDNS_7246548160561 $T=285215 135035 0 0 $X=284245 $Y=134895
X331 2 VIA1_C_CDNS_7246548160561 $T=285215 153835 0 0 $X=284245 $Y=153695
X332 30 VIA1_C_CDNS_7246548160561 $T=293585 115455 0 0 $X=292615 $Y=115315
X333 2 VIA1_C_CDNS_7246548160561 $T=296455 78635 0 0 $X=295485 $Y=78495
X334 2 VIA1_C_CDNS_7246548160561 $T=296455 97435 0 0 $X=295485 $Y=97295
X335 2 VIA1_C_CDNS_7246548160561 $T=296455 116235 0 0 $X=295485 $Y=116095
X336 2 VIA1_C_CDNS_7246548160561 $T=296455 135035 0 0 $X=295485 $Y=134895
X337 2 VIA1_C_CDNS_7246548160561 $T=296455 153835 0 0 $X=295485 $Y=153695
X338 28 VIA1_C_CDNS_7246548160561 $T=304825 113115 0 0 $X=303855 $Y=112975
X339 2 VIA1_C_CDNS_7246548160561 $T=307695 78635 0 0 $X=306725 $Y=78495
X340 2 VIA1_C_CDNS_7246548160561 $T=307695 97435 0 0 $X=306725 $Y=97295
X341 2 VIA1_C_CDNS_7246548160561 $T=307695 116235 0 0 $X=306725 $Y=116095
X342 2 VIA1_C_CDNS_7246548160561 $T=307695 135035 0 0 $X=306725 $Y=134895
X343 2 VIA1_C_CDNS_7246548160561 $T=307695 153835 0 0 $X=306725 $Y=153695
X344 27 VIA1_C_CDNS_7246548160561 $T=316065 113895 0 0 $X=315095 $Y=113755
X345 2 VIA1_C_CDNS_7246548160561 $T=318315 78635 0 0 $X=317345 $Y=78495
X346 2 VIA1_C_CDNS_7246548160561 $T=318935 97435 0 0 $X=317965 $Y=97295
X347 2 VIA1_C_CDNS_7246548160561 $T=318935 116235 0 0 $X=317965 $Y=116095
X348 2 VIA1_C_CDNS_7246548160561 $T=318935 135035 0 0 $X=317965 $Y=134895
X349 2 VIA1_C_CDNS_7246548160561 $T=318935 153835 0 0 $X=317965 $Y=153695
X350 26 VIA1_C_CDNS_7246548160561 $T=327305 114675 0 0 $X=326335 $Y=114535
X351 2 VIA1_C_CDNS_7246548160561 $T=329555 78635 0 0 $X=328585 $Y=78495
X352 2 VIA1_C_CDNS_7246548160561 $T=330175 97435 0 0 $X=329205 $Y=97295
X353 2 VIA1_C_CDNS_7246548160561 $T=330175 116235 0 0 $X=329205 $Y=116095
X354 2 VIA1_C_CDNS_7246548160561 $T=330175 135035 0 0 $X=329205 $Y=134895
X355 2 VIA1_C_CDNS_7246548160561 $T=330175 153835 0 0 $X=329205 $Y=153695
X356 26 VIA1_C_CDNS_7246548160561 $T=338545 114675 0 0 $X=337575 $Y=114535
X357 2 VIA1_C_CDNS_7246548160561 $T=340795 78635 0 0 $X=339825 $Y=78495
X358 2 VIA1_C_CDNS_7246548160561 $T=341415 97435 0 0 $X=340445 $Y=97295
X359 2 VIA1_C_CDNS_7246548160561 $T=341415 116235 0 0 $X=340445 $Y=116095
X360 2 VIA1_C_CDNS_7246548160561 $T=341415 135035 0 0 $X=340445 $Y=134895
X361 2 VIA1_C_CDNS_7246548160561 $T=341415 153835 0 0 $X=340445 $Y=153695
X362 26 VIA1_C_CDNS_7246548160561 $T=349785 114675 0 0 $X=348815 $Y=114535
X363 2 VIA1_C_CDNS_7246548160561 $T=352035 78635 0 0 $X=351065 $Y=78495
X364 2 VIA1_C_CDNS_7246548160561 $T=352655 97435 0 0 $X=351685 $Y=97295
X365 2 VIA1_C_CDNS_7246548160561 $T=352655 116235 0 0 $X=351685 $Y=116095
X366 2 VIA1_C_CDNS_7246548160561 $T=352655 135035 0 0 $X=351685 $Y=134895
X367 2 VIA1_C_CDNS_7246548160561 $T=352655 153835 0 0 $X=351685 $Y=153695
X368 26 VIA1_C_CDNS_7246548160561 $T=361025 114675 0 0 $X=360055 $Y=114535
X369 2 VIA1_C_CDNS_7246548160561 $T=363275 78635 0 0 $X=362305 $Y=78495
X370 2 VIA1_C_CDNS_7246548160561 $T=363845 97435 0 0 $X=362875 $Y=97295
X371 2 VIA1_C_CDNS_7246548160561 $T=363845 116235 0 0 $X=362875 $Y=116095
X372 2 VIA1_C_CDNS_7246548160561 $T=363845 135035 0 0 $X=362875 $Y=134895
X373 2 VIA1_C_CDNS_7246548160561 $T=363845 153835 0 0 $X=362875 $Y=153695
X374 2 VIA1_C_CDNS_7246548160562 $T=205165 59835 0 0 $X=204245 $Y=59645
X375 2 VIA1_C_CDNS_7246548160562 $T=205165 78635 0 0 $X=204245 $Y=78445
X376 2 VIA1_C_CDNS_7246548160562 $T=205165 97435 0 0 $X=204245 $Y=97245
X377 2 VIA1_C_CDNS_7246548160562 $T=205165 116235 0 0 $X=204245 $Y=116045
X378 2 VIA1_C_CDNS_7246548160562 $T=205165 135035 0 0 $X=204245 $Y=134845
X379 2 VIA1_C_CDNS_7246548160562 $T=205165 153835 0 0 $X=204245 $Y=153645
X380 2 VIA1_C_CDNS_7246548160562 $T=205165 172635 0 0 $X=204245 $Y=172445
X381 2 VIA1_C_CDNS_7246548160562 $T=205165 177475 0 0 $X=204245 $Y=177285
X382 2 VIA1_C_CDNS_7246548160562 $T=210435 48755 0 0 $X=209515 $Y=48565
X383 2 VIA1_C_CDNS_7246548160562 $T=210435 59835 0 0 $X=209515 $Y=59645
X384 2 VIA1_C_CDNS_7246548160562 $T=210435 78635 0 0 $X=209515 $Y=78445
X385 2 VIA1_C_CDNS_7246548160562 $T=210435 97435 0 0 $X=209515 $Y=97245
X386 2 VIA1_C_CDNS_7246548160562 $T=210435 116235 0 0 $X=209515 $Y=116045
X387 2 VIA1_C_CDNS_7246548160562 $T=210435 135035 0 0 $X=209515 $Y=134845
X388 2 VIA1_C_CDNS_7246548160562 $T=210435 153835 0 0 $X=209515 $Y=153645
X389 2 VIA1_C_CDNS_7246548160562 $T=210435 172635 0 0 $X=209515 $Y=172445
X390 2 VIA1_C_CDNS_7246548160562 $T=214955 59835 0 0 $X=214035 $Y=59645
X391 2 VIA1_C_CDNS_7246548160562 $T=214955 78635 0 0 $X=214035 $Y=78445
X392 2 VIA1_C_CDNS_7246548160562 $T=214955 97435 0 0 $X=214035 $Y=97245
X393 2 VIA1_C_CDNS_7246548160562 $T=214955 135035 0 0 $X=214035 $Y=134845
X394 2 VIA1_C_CDNS_7246548160562 $T=214955 153835 0 0 $X=214035 $Y=153645
X395 2 VIA1_C_CDNS_7246548160562 $T=214955 172635 0 0 $X=214035 $Y=172445
X396 2 VIA1_C_CDNS_7246548160562 $T=214955 177475 0 0 $X=214035 $Y=177285
X397 2 VIA1_C_CDNS_7246548160562 $T=217155 59835 0 0 $X=216235 $Y=59645
X398 2 VIA1_C_CDNS_7246548160562 $T=217155 172635 0 0 $X=216235 $Y=172445
X399 2 VIA1_C_CDNS_7246548160562 $T=217155 177475 0 0 $X=216235 $Y=177285
X400 2 VIA1_C_CDNS_7246548160562 $T=221675 48755 0 0 $X=220755 $Y=48565
X401 17 VIA1_C_CDNS_7246548160562 $T=221675 54375 0 0 $X=220755 $Y=54185
X402 17 VIA1_C_CDNS_7246548160562 $T=221675 73175 0 0 $X=220755 $Y=72985
X403 17 VIA1_C_CDNS_7246548160562 $T=221675 91975 0 0 $X=220755 $Y=91785
X404 17 VIA1_C_CDNS_7246548160562 $T=221675 110775 0 0 $X=220755 $Y=110585
X405 17 VIA1_C_CDNS_7246548160562 $T=221675 129575 0 0 $X=220755 $Y=129385
X406 17 VIA1_C_CDNS_7246548160562 $T=221675 148375 0 0 $X=220755 $Y=148185
X407 2 VIA1_C_CDNS_7246548160562 $T=221675 172635 0 0 $X=220755 $Y=172445
X408 2 VIA1_C_CDNS_7246548160562 $T=226195 59835 0 0 $X=225275 $Y=59645
X409 26 VIA1_C_CDNS_7246548160562 $T=226195 77075 0 0 $X=225275 $Y=76885
X410 26 VIA1_C_CDNS_7246548160562 $T=226195 95875 0 0 $X=225275 $Y=95685
X411 26 VIA1_C_CDNS_7246548160562 $T=226195 133475 0 0 $X=225275 $Y=133285
X412 26 VIA1_C_CDNS_7246548160562 $T=226195 152275 0 0 $X=225275 $Y=152085
X413 26 VIA1_C_CDNS_7246548160562 $T=226195 171075 0 0 $X=225275 $Y=170885
X414 2 VIA1_C_CDNS_7246548160562 $T=226195 177475 0 0 $X=225275 $Y=177285
X415 2 VIA1_C_CDNS_7246548160562 $T=228395 59835 0 0 $X=227475 $Y=59645
X416 2 VIA1_C_CDNS_7246548160562 $T=228395 177475 0 0 $X=227475 $Y=177285
X417 2 VIA1_C_CDNS_7246548160562 $T=228965 172635 0 0 $X=228045 $Y=172445
X418 2 VIA1_C_CDNS_7246548160562 $T=232915 48755 0 0 $X=231995 $Y=48565
X419 17 VIA1_C_CDNS_7246548160562 $T=232915 54375 0 0 $X=231995 $Y=54185
X420 17 VIA1_C_CDNS_7246548160562 $T=232915 73175 0 0 $X=231995 $Y=72985
X421 17 VIA1_C_CDNS_7246548160562 $T=232915 91975 0 0 $X=231995 $Y=91785
X422 17 VIA1_C_CDNS_7246548160562 $T=232915 110775 0 0 $X=231995 $Y=110585
X423 17 VIA1_C_CDNS_7246548160562 $T=232915 129575 0 0 $X=231995 $Y=129385
X424 17 VIA1_C_CDNS_7246548160562 $T=232915 148375 0 0 $X=231995 $Y=148185
X425 2 VIA1_C_CDNS_7246548160562 $T=232915 172635 0 0 $X=231995 $Y=172445
X426 2 VIA1_C_CDNS_7246548160562 $T=237435 59835 0 0 $X=236515 $Y=59645
X427 27 VIA1_C_CDNS_7246548160562 $T=237435 76295 0 0 $X=236515 $Y=76105
X428 27 VIA1_C_CDNS_7246548160562 $T=237435 95095 0 0 $X=236515 $Y=94905
X429 27 VIA1_C_CDNS_7246548160562 $T=237435 132695 0 0 $X=236515 $Y=132505
X430 27 VIA1_C_CDNS_7246548160562 $T=237435 151495 0 0 $X=236515 $Y=151305
X431 26 VIA1_C_CDNS_7246548160562 $T=237435 171075 0 0 $X=236515 $Y=170885
X432 2 VIA1_C_CDNS_7246548160562 $T=237435 177475 0 0 $X=236515 $Y=177285
X433 2 VIA1_C_CDNS_7246548160562 $T=239635 59835 0 0 $X=238715 $Y=59645
X434 2 VIA1_C_CDNS_7246548160562 $T=239635 177475 0 0 $X=238715 $Y=177285
X435 2 VIA1_C_CDNS_7246548160562 $T=240205 172635 0 0 $X=239285 $Y=172445
X436 2 VIA1_C_CDNS_7246548160562 $T=244155 48755 0 0 $X=243235 $Y=48565
X437 17 VIA1_C_CDNS_7246548160562 $T=244155 54375 0 0 $X=243235 $Y=54185
X438 17 VIA1_C_CDNS_7246548160562 $T=244155 73175 0 0 $X=243235 $Y=72985
X439 17 VIA1_C_CDNS_7246548160562 $T=244155 91975 0 0 $X=243235 $Y=91785
X440 17 VIA1_C_CDNS_7246548160562 $T=244155 110775 0 0 $X=243235 $Y=110585
X441 17 VIA1_C_CDNS_7246548160562 $T=244155 129575 0 0 $X=243235 $Y=129385
X442 17 VIA1_C_CDNS_7246548160562 $T=244155 148375 0 0 $X=243235 $Y=148185
X443 2 VIA1_C_CDNS_7246548160562 $T=244155 172635 0 0 $X=243235 $Y=172445
X444 2 VIA1_C_CDNS_7246548160562 $T=248675 59835 0 0 $X=247755 $Y=59645
X445 27 VIA1_C_CDNS_7246548160562 $T=248675 76295 0 0 $X=247755 $Y=76105
X446 28 VIA1_C_CDNS_7246548160562 $T=248675 94315 0 0 $X=247755 $Y=94125
X447 28 VIA1_C_CDNS_7246548160562 $T=248675 131915 0 0 $X=247755 $Y=131725
X448 28 VIA1_C_CDNS_7246548160562 $T=248675 150715 0 0 $X=247755 $Y=150525
X449 26 VIA1_C_CDNS_7246548160562 $T=248675 171075 0 0 $X=247755 $Y=170885
X450 2 VIA1_C_CDNS_7246548160562 $T=248675 177475 0 0 $X=247755 $Y=177285
X451 2 VIA1_C_CDNS_7246548160562 $T=250875 59835 0 0 $X=249955 $Y=59645
X452 2 VIA1_C_CDNS_7246548160562 $T=250875 177475 0 0 $X=249955 $Y=177285
X453 2 VIA1_C_CDNS_7246548160562 $T=251445 172635 0 0 $X=250525 $Y=172445
X454 2 VIA1_C_CDNS_7246548160562 $T=255395 48755 0 0 $X=254475 $Y=48565
X455 17 VIA1_C_CDNS_7246548160562 $T=255395 54375 0 0 $X=254475 $Y=54185
X456 17 VIA1_C_CDNS_7246548160562 $T=255395 73175 0 0 $X=254475 $Y=72985
X457 17 VIA1_C_CDNS_7246548160562 $T=255395 91975 0 0 $X=254475 $Y=91785
X458 17 VIA1_C_CDNS_7246548160562 $T=255395 110775 0 0 $X=254475 $Y=110585
X459 17 VIA1_C_CDNS_7246548160562 $T=255395 129575 0 0 $X=254475 $Y=129385
X460 17 VIA1_C_CDNS_7246548160562 $T=255395 148375 0 0 $X=254475 $Y=148185
X461 2 VIA1_C_CDNS_7246548160562 $T=255395 172635 0 0 $X=254475 $Y=172445
X462 2 VIA1_C_CDNS_7246548160562 $T=259915 59835 0 0 $X=258995 $Y=59645
X463 27 VIA1_C_CDNS_7246548160562 $T=259915 76295 0 0 $X=258995 $Y=76105
X464 30 VIA1_C_CDNS_7246548160562 $T=259915 96655 0 0 $X=258995 $Y=96465
X465 30 VIA1_C_CDNS_7246548160562 $T=259915 134255 0 0 $X=258995 $Y=134065
X466 30 VIA1_C_CDNS_7246548160562 $T=259915 153055 0 0 $X=258995 $Y=152865
X467 26 VIA1_C_CDNS_7246548160562 $T=259915 171075 0 0 $X=258995 $Y=170885
X468 2 VIA1_C_CDNS_7246548160562 $T=259915 177475 0 0 $X=258995 $Y=177285
X469 2 VIA1_C_CDNS_7246548160562 $T=262115 59835 0 0 $X=261195 $Y=59645
X470 2 VIA1_C_CDNS_7246548160562 $T=262115 177475 0 0 $X=261195 $Y=177285
X471 2 VIA1_C_CDNS_7246548160562 $T=262685 172635 0 0 $X=261765 $Y=172445
X472 2 VIA1_C_CDNS_7246548160562 $T=266635 48755 0 0 $X=265715 $Y=48565
X473 17 VIA1_C_CDNS_7246548160562 $T=266635 54375 0 0 $X=265715 $Y=54185
X474 17 VIA1_C_CDNS_7246548160562 $T=266635 73175 0 0 $X=265715 $Y=72985
X475 17 VIA1_C_CDNS_7246548160562 $T=266635 91975 0 0 $X=265715 $Y=91785
X476 17 VIA1_C_CDNS_7246548160562 $T=266635 110775 0 0 $X=265715 $Y=110585
X477 17 VIA1_C_CDNS_7246548160562 $T=266635 129575 0 0 $X=265715 $Y=129385
X478 17 VIA1_C_CDNS_7246548160562 $T=266635 148375 0 0 $X=265715 $Y=148185
X479 2 VIA1_C_CDNS_7246548160562 $T=266635 172635 0 0 $X=265715 $Y=172445
X480 2 VIA1_C_CDNS_7246548160562 $T=271155 59835 0 0 $X=270235 $Y=59645
X481 27 VIA1_C_CDNS_7246548160562 $T=271155 76295 0 0 $X=270235 $Y=76105
X482 31 VIA1_C_CDNS_7246548160562 $T=271155 93535 0 0 $X=270235 $Y=93345
X483 29 VIA1_C_CDNS_7246548160562 $T=271155 130355 0 0 $X=270235 $Y=130165
X484 31 VIA1_C_CDNS_7246548160562 $T=271155 149935 0 0 $X=270235 $Y=149745
X485 26 VIA1_C_CDNS_7246548160562 $T=271155 171075 0 0 $X=270235 $Y=170885
X486 2 VIA1_C_CDNS_7246548160562 $T=271155 177475 0 0 $X=270235 $Y=177285
X487 2 VIA1_C_CDNS_7246548160562 $T=273355 59835 0 0 $X=272435 $Y=59645
X488 2 VIA1_C_CDNS_7246548160562 $T=273355 177475 0 0 $X=272435 $Y=177285
X489 2 VIA1_C_CDNS_7246548160562 $T=273925 172635 0 0 $X=273005 $Y=172445
X490 2 VIA1_C_CDNS_7246548160562 $T=277875 48755 0 0 $X=276955 $Y=48565
X491 17 VIA1_C_CDNS_7246548160562 $T=277875 54375 0 0 $X=276955 $Y=54185
X492 17 VIA1_C_CDNS_7246548160562 $T=277875 73175 0 0 $X=276955 $Y=72985
X493 17 VIA1_C_CDNS_7246548160562 $T=277875 91975 0 0 $X=276955 $Y=91785
X494 17 VIA1_C_CDNS_7246548160562 $T=277875 110775 0 0 $X=276955 $Y=110585
X495 17 VIA1_C_CDNS_7246548160562 $T=277875 129575 0 0 $X=276955 $Y=129385
X496 17 VIA1_C_CDNS_7246548160562 $T=277875 148375 0 0 $X=276955 $Y=148185
X497 2 VIA1_C_CDNS_7246548160562 $T=277875 172635 0 0 $X=276955 $Y=172445
X498 2 VIA1_C_CDNS_7246548160562 $T=282395 59835 0 0 $X=281475 $Y=59645
X499 30 VIA1_C_CDNS_7246548160562 $T=282395 77855 0 0 $X=281475 $Y=77665
X500 31 VIA1_C_CDNS_7246548160562 $T=282395 93535 0 0 $X=281475 $Y=93345
X501 30 VIA1_C_CDNS_7246548160562 $T=282395 134255 0 0 $X=281475 $Y=134065
X502 31 VIA1_C_CDNS_7246548160562 $T=282395 149935 0 0 $X=281475 $Y=149745
X503 27 VIA1_C_CDNS_7246548160562 $T=282395 170295 0 0 $X=281475 $Y=170105
X504 2 VIA1_C_CDNS_7246548160562 $T=282395 177475 0 0 $X=281475 $Y=177285
X505 2 VIA1_C_CDNS_7246548160562 $T=284595 59835 0 0 $X=283675 $Y=59645
X506 2 VIA1_C_CDNS_7246548160562 $T=284595 177475 0 0 $X=283675 $Y=177285
X507 2 VIA1_C_CDNS_7246548160562 $T=285165 172635 0 0 $X=284245 $Y=172445
X508 2 VIA1_C_CDNS_7246548160562 $T=289115 48755 0 0 $X=288195 $Y=48565
X509 17 VIA1_C_CDNS_7246548160562 $T=289115 54375 0 0 $X=288195 $Y=54185
X510 17 VIA1_C_CDNS_7246548160562 $T=289115 73175 0 0 $X=288195 $Y=72985
X511 17 VIA1_C_CDNS_7246548160562 $T=289115 91975 0 0 $X=288195 $Y=91785
X512 17 VIA1_C_CDNS_7246548160562 $T=289115 110775 0 0 $X=288195 $Y=110585
X513 17 VIA1_C_CDNS_7246548160562 $T=289115 129575 0 0 $X=288195 $Y=129385
X514 17 VIA1_C_CDNS_7246548160562 $T=289115 148375 0 0 $X=288195 $Y=148185
X515 2 VIA1_C_CDNS_7246548160562 $T=289115 172635 0 0 $X=288195 $Y=172445
X516 2 VIA1_C_CDNS_7246548160562 $T=293635 59835 0 0 $X=292715 $Y=59645
X517 26 VIA1_C_CDNS_7246548160562 $T=293635 77075 0 0 $X=292715 $Y=76885
X518 30 VIA1_C_CDNS_7246548160562 $T=293635 96655 0 0 $X=292715 $Y=96465
X519 28 VIA1_C_CDNS_7246548160562 $T=293635 131915 0 0 $X=292715 $Y=131725
X520 30 VIA1_C_CDNS_7246548160562 $T=293635 153055 0 0 $X=292715 $Y=152865
X521 27 VIA1_C_CDNS_7246548160562 $T=293635 170295 0 0 $X=292715 $Y=170105
X522 2 VIA1_C_CDNS_7246548160562 $T=293635 177475 0 0 $X=292715 $Y=177285
X523 2 VIA1_C_CDNS_7246548160562 $T=295835 59835 0 0 $X=294915 $Y=59645
X524 2 VIA1_C_CDNS_7246548160562 $T=295835 177475 0 0 $X=294915 $Y=177285
X525 2 VIA1_C_CDNS_7246548160562 $T=296405 172635 0 0 $X=295485 $Y=172445
X526 2 VIA1_C_CDNS_7246548160562 $T=300355 48755 0 0 $X=299435 $Y=48565
X527 17 VIA1_C_CDNS_7246548160562 $T=300355 54375 0 0 $X=299435 $Y=54185
X528 17 VIA1_C_CDNS_7246548160562 $T=300355 73175 0 0 $X=299435 $Y=72985
X529 17 VIA1_C_CDNS_7246548160562 $T=300355 91975 0 0 $X=299435 $Y=91785
X530 17 VIA1_C_CDNS_7246548160562 $T=300355 110775 0 0 $X=299435 $Y=110585
X531 17 VIA1_C_CDNS_7246548160562 $T=300355 129575 0 0 $X=299435 $Y=129385
X532 17 VIA1_C_CDNS_7246548160562 $T=300355 148375 0 0 $X=299435 $Y=148185
X533 2 VIA1_C_CDNS_7246548160562 $T=300355 172635 0 0 $X=299435 $Y=172445
X534 2 VIA1_C_CDNS_7246548160562 $T=304875 59835 0 0 $X=303955 $Y=59645
X535 26 VIA1_C_CDNS_7246548160562 $T=304875 77075 0 0 $X=303955 $Y=76885
X536 28 VIA1_C_CDNS_7246548160562 $T=304875 94315 0 0 $X=303955 $Y=94125
X537 27 VIA1_C_CDNS_7246548160562 $T=304875 132695 0 0 $X=303955 $Y=132505
X538 28 VIA1_C_CDNS_7246548160562 $T=304875 150715 0 0 $X=303955 $Y=150525
X539 27 VIA1_C_CDNS_7246548160562 $T=304875 170295 0 0 $X=303955 $Y=170105
X540 2 VIA1_C_CDNS_7246548160562 $T=304875 177475 0 0 $X=303955 $Y=177285
X541 2 VIA1_C_CDNS_7246548160562 $T=307075 59835 0 0 $X=306155 $Y=59645
X542 2 VIA1_C_CDNS_7246548160562 $T=307075 177475 0 0 $X=306155 $Y=177285
X543 2 VIA1_C_CDNS_7246548160562 $T=307645 172635 0 0 $X=306725 $Y=172445
X544 2 VIA1_C_CDNS_7246548160562 $T=311595 48755 0 0 $X=310675 $Y=48565
X545 2 VIA1_C_CDNS_7246548160562 $T=311595 59835 0 0 $X=310675 $Y=59645
X546 17 VIA1_C_CDNS_7246548160562 $T=311595 73175 0 0 $X=310675 $Y=72985
X547 17 VIA1_C_CDNS_7246548160562 $T=311595 91975 0 0 $X=310675 $Y=91785
X548 17 VIA1_C_CDNS_7246548160562 $T=311595 110775 0 0 $X=310675 $Y=110585
X549 17 VIA1_C_CDNS_7246548160562 $T=311595 129575 0 0 $X=310675 $Y=129385
X550 17 VIA1_C_CDNS_7246548160562 $T=311595 148375 0 0 $X=310675 $Y=148185
X551 2 VIA1_C_CDNS_7246548160562 $T=311595 172635 0 0 $X=310675 $Y=172445
X552 2 VIA1_C_CDNS_7246548160562 $T=316115 59835 0 0 $X=315195 $Y=59645
X553 2 VIA1_C_CDNS_7246548160562 $T=316115 78635 0 0 $X=315195 $Y=78445
X554 27 VIA1_C_CDNS_7246548160562 $T=316115 95095 0 0 $X=315195 $Y=94905
X555 27 VIA1_C_CDNS_7246548160562 $T=316115 132695 0 0 $X=315195 $Y=132505
X556 27 VIA1_C_CDNS_7246548160562 $T=316115 151495 0 0 $X=315195 $Y=151305
X557 30 VIA1_C_CDNS_7246548160562 $T=316115 171855 0 0 $X=315195 $Y=171665
X558 2 VIA1_C_CDNS_7246548160562 $T=316115 177475 0 0 $X=315195 $Y=177285
X559 2 VIA1_C_CDNS_7246548160562 $T=318315 59835 0 0 $X=317395 $Y=59645
X560 2 VIA1_C_CDNS_7246548160562 $T=318315 177475 0 0 $X=317395 $Y=177285
X561 2 VIA1_C_CDNS_7246548160562 $T=318885 172635 0 0 $X=317965 $Y=172445
X562 2 VIA1_C_CDNS_7246548160562 $T=322835 48755 0 0 $X=321915 $Y=48565
X563 2 VIA1_C_CDNS_7246548160562 $T=322835 59835 0 0 $X=321915 $Y=59645
X564 17 VIA1_C_CDNS_7246548160562 $T=322835 73175 0 0 $X=321915 $Y=72985
X565 17 VIA1_C_CDNS_7246548160562 $T=322835 91975 0 0 $X=321915 $Y=91785
X566 17 VIA1_C_CDNS_7246548160562 $T=322835 110775 0 0 $X=321915 $Y=110585
X567 17 VIA1_C_CDNS_7246548160562 $T=322835 129575 0 0 $X=321915 $Y=129385
X568 17 VIA1_C_CDNS_7246548160562 $T=322835 148375 0 0 $X=321915 $Y=148185
X569 2 VIA1_C_CDNS_7246548160562 $T=322835 172635 0 0 $X=321915 $Y=172445
X570 2 VIA1_C_CDNS_7246548160562 $T=327355 59835 0 0 $X=326435 $Y=59645
X571 2 VIA1_C_CDNS_7246548160562 $T=327355 78635 0 0 $X=326435 $Y=78445
X572 26 VIA1_C_CDNS_7246548160562 $T=327355 95875 0 0 $X=326435 $Y=95685
X573 26 VIA1_C_CDNS_7246548160562 $T=327355 133475 0 0 $X=326435 $Y=133285
X574 26 VIA1_C_CDNS_7246548160562 $T=327355 152275 0 0 $X=326435 $Y=152085
X575 26 VIA1_C_CDNS_7246548160562 $T=327355 171075 0 0 $X=326435 $Y=170885
X576 2 VIA1_C_CDNS_7246548160562 $T=327355 177475 0 0 $X=326435 $Y=177285
X577 2 VIA1_C_CDNS_7246548160562 $T=329555 59835 0 0 $X=328635 $Y=59645
X578 2 VIA1_C_CDNS_7246548160562 $T=329555 177475 0 0 $X=328635 $Y=177285
X579 2 VIA1_C_CDNS_7246548160562 $T=330125 172635 0 0 $X=329205 $Y=172445
X580 2 VIA1_C_CDNS_7246548160562 $T=334075 48755 0 0 $X=333155 $Y=48565
X581 2 VIA1_C_CDNS_7246548160562 $T=334075 59835 0 0 $X=333155 $Y=59645
X582 17 VIA1_C_CDNS_7246548160562 $T=334075 73175 0 0 $X=333155 $Y=72985
X583 17 VIA1_C_CDNS_7246548160562 $T=334075 91975 0 0 $X=333155 $Y=91785
X584 17 VIA1_C_CDNS_7246548160562 $T=334075 110775 0 0 $X=333155 $Y=110585
X585 17 VIA1_C_CDNS_7246548160562 $T=334075 129575 0 0 $X=333155 $Y=129385
X586 17 VIA1_C_CDNS_7246548160562 $T=334075 148375 0 0 $X=333155 $Y=148185
X587 2 VIA1_C_CDNS_7246548160562 $T=334075 172635 0 0 $X=333155 $Y=172445
X588 2 VIA1_C_CDNS_7246548160562 $T=338595 59835 0 0 $X=337675 $Y=59645
X589 2 VIA1_C_CDNS_7246548160562 $T=338595 78635 0 0 $X=337675 $Y=78445
X590 26 VIA1_C_CDNS_7246548160562 $T=338595 95875 0 0 $X=337675 $Y=95685
X591 26 VIA1_C_CDNS_7246548160562 $T=338595 133475 0 0 $X=337675 $Y=133285
X592 26 VIA1_C_CDNS_7246548160562 $T=338595 152275 0 0 $X=337675 $Y=152085
X593 26 VIA1_C_CDNS_7246548160562 $T=338595 171075 0 0 $X=337675 $Y=170885
X594 2 VIA1_C_CDNS_7246548160562 $T=338595 177475 0 0 $X=337675 $Y=177285
X595 2 VIA1_C_CDNS_7246548160562 $T=340795 59835 0 0 $X=339875 $Y=59645
X596 2 VIA1_C_CDNS_7246548160562 $T=340795 177475 0 0 $X=339875 $Y=177285
X597 2 VIA1_C_CDNS_7246548160562 $T=341365 172635 0 0 $X=340445 $Y=172445
X598 2 VIA1_C_CDNS_7246548160562 $T=345315 48755 0 0 $X=344395 $Y=48565
X599 2 VIA1_C_CDNS_7246548160562 $T=345315 59835 0 0 $X=344395 $Y=59645
X600 17 VIA1_C_CDNS_7246548160562 $T=345315 73175 0 0 $X=344395 $Y=72985
X601 17 VIA1_C_CDNS_7246548160562 $T=345315 91975 0 0 $X=344395 $Y=91785
X602 17 VIA1_C_CDNS_7246548160562 $T=345315 110775 0 0 $X=344395 $Y=110585
X603 17 VIA1_C_CDNS_7246548160562 $T=345315 129575 0 0 $X=344395 $Y=129385
X604 17 VIA1_C_CDNS_7246548160562 $T=345315 148375 0 0 $X=344395 $Y=148185
X605 2 VIA1_C_CDNS_7246548160562 $T=345315 172635 0 0 $X=344395 $Y=172445
X606 2 VIA1_C_CDNS_7246548160562 $T=349835 59835 0 0 $X=348915 $Y=59645
X607 2 VIA1_C_CDNS_7246548160562 $T=349835 78635 0 0 $X=348915 $Y=78445
X608 26 VIA1_C_CDNS_7246548160562 $T=349835 95875 0 0 $X=348915 $Y=95685
X609 26 VIA1_C_CDNS_7246548160562 $T=349835 133475 0 0 $X=348915 $Y=133285
X610 26 VIA1_C_CDNS_7246548160562 $T=349835 152275 0 0 $X=348915 $Y=152085
X611 26 VIA1_C_CDNS_7246548160562 $T=349835 171075 0 0 $X=348915 $Y=170885
X612 2 VIA1_C_CDNS_7246548160562 $T=349835 177475 0 0 $X=348915 $Y=177285
X613 2 VIA1_C_CDNS_7246548160562 $T=352035 59835 0 0 $X=351115 $Y=59645
X614 2 VIA1_C_CDNS_7246548160562 $T=352035 177475 0 0 $X=351115 $Y=177285
X615 2 VIA1_C_CDNS_7246548160562 $T=352605 172635 0 0 $X=351685 $Y=172445
X616 2 VIA1_C_CDNS_7246548160562 $T=356555 48755 0 0 $X=355635 $Y=48565
X617 2 VIA1_C_CDNS_7246548160562 $T=356555 59835 0 0 $X=355635 $Y=59645
X618 17 VIA1_C_CDNS_7246548160562 $T=356555 73175 0 0 $X=355635 $Y=72985
X619 17 VIA1_C_CDNS_7246548160562 $T=356555 91975 0 0 $X=355635 $Y=91785
X620 17 VIA1_C_CDNS_7246548160562 $T=356555 110775 0 0 $X=355635 $Y=110585
X621 17 VIA1_C_CDNS_7246548160562 $T=356555 129575 0 0 $X=355635 $Y=129385
X622 17 VIA1_C_CDNS_7246548160562 $T=356555 148375 0 0 $X=355635 $Y=148185
X623 2 VIA1_C_CDNS_7246548160562 $T=356555 172635 0 0 $X=355635 $Y=172445
X624 2 VIA1_C_CDNS_7246548160562 $T=361075 59835 0 0 $X=360155 $Y=59645
X625 2 VIA1_C_CDNS_7246548160562 $T=361075 78635 0 0 $X=360155 $Y=78445
X626 26 VIA1_C_CDNS_7246548160562 $T=361075 95875 0 0 $X=360155 $Y=95685
X627 26 VIA1_C_CDNS_7246548160562 $T=361075 133475 0 0 $X=360155 $Y=133285
X628 26 VIA1_C_CDNS_7246548160562 $T=361075 152275 0 0 $X=360155 $Y=152085
X629 26 VIA1_C_CDNS_7246548160562 $T=361075 171075 0 0 $X=360155 $Y=170885
X630 2 VIA1_C_CDNS_7246548160562 $T=361075 177475 0 0 $X=360155 $Y=177285
X631 2 VIA1_C_CDNS_7246548160562 $T=363275 59835 0 0 $X=362355 $Y=59645
X632 2 VIA1_C_CDNS_7246548160562 $T=363275 177475 0 0 $X=362355 $Y=177285
X633 2 VIA1_C_CDNS_7246548160562 $T=363845 172635 0 0 $X=362925 $Y=172445
X634 2 VIA1_C_CDNS_7246548160562 $T=367795 48755 0 0 $X=366875 $Y=48565
X635 2 VIA1_C_CDNS_7246548160562 $T=367795 59835 0 0 $X=366875 $Y=59645
X636 2 VIA1_C_CDNS_7246548160562 $T=367795 78635 0 0 $X=366875 $Y=78445
X637 2 VIA1_C_CDNS_7246548160562 $T=367795 97435 0 0 $X=366875 $Y=97245
X638 2 VIA1_C_CDNS_7246548160562 $T=367795 116235 0 0 $X=366875 $Y=116045
X639 2 VIA1_C_CDNS_7246548160562 $T=367795 135035 0 0 $X=366875 $Y=134845
X640 2 VIA1_C_CDNS_7246548160562 $T=367795 153835 0 0 $X=366875 $Y=153645
X641 2 VIA1_C_CDNS_7246548160562 $T=367795 172635 0 0 $X=366875 $Y=172445
X642 2 VIA1_C_CDNS_7246548160562 $T=373065 59835 0 0 $X=372145 $Y=59645
X643 2 VIA1_C_CDNS_7246548160562 $T=373065 78635 0 0 $X=372145 $Y=78445
X644 2 VIA1_C_CDNS_7246548160562 $T=373065 97435 0 0 $X=372145 $Y=97245
X645 2 VIA1_C_CDNS_7246548160562 $T=373065 116235 0 0 $X=372145 $Y=116045
X646 2 VIA1_C_CDNS_7246548160562 $T=373065 135035 0 0 $X=372145 $Y=134845
X647 2 VIA1_C_CDNS_7246548160562 $T=373065 153835 0 0 $X=372145 $Y=153645
X648 2 VIA1_C_CDNS_7246548160562 $T=373065 172635 0 0 $X=372145 $Y=172445
X649 2 VIA1_C_CDNS_7246548160562 $T=373065 177475 0 0 $X=372145 $Y=177285
X650 24 VIA2_C_CDNS_7246548160563 $T=184405 53595 0 0 $X=183485 $Y=53405
X651 24 VIA2_C_CDNS_7246548160563 $T=184405 72395 0 0 $X=183485 $Y=72205
X652 24 VIA2_C_CDNS_7246548160563 $T=184405 91195 0 0 $X=183485 $Y=91005
X653 24 VIA2_C_CDNS_7246548160563 $T=184405 109995 0 0 $X=183485 $Y=109805
X654 24 VIA2_C_CDNS_7246548160563 $T=184405 128795 0 0 $X=183485 $Y=128605
X655 24 VIA2_C_CDNS_7246548160563 $T=184405 147595 0 0 $X=183485 $Y=147405
X656 24 VIA2_C_CDNS_7246548160563 $T=184405 166395 0 0 $X=183485 $Y=166205
X657 17 VIA2_C_CDNS_7246548160563 $T=186685 54375 0 0 $X=185765 $Y=54185
X658 17 VIA2_C_CDNS_7246548160563 $T=186685 73175 0 0 $X=185765 $Y=72985
X659 17 VIA2_C_CDNS_7246548160563 $T=186685 91975 0 0 $X=185765 $Y=91785
X660 17 VIA2_C_CDNS_7246548160563 $T=186685 110775 0 0 $X=185765 $Y=110585
X661 17 VIA2_C_CDNS_7246548160563 $T=186685 129575 0 0 $X=185765 $Y=129385
X662 17 VIA2_C_CDNS_7246548160563 $T=186685 148375 0 0 $X=185765 $Y=148185
X663 17 VIA2_C_CDNS_7246548160563 $T=186685 167175 0 0 $X=185765 $Y=166985
X664 29 VIA2_C_CDNS_7246548160563 $T=188965 55155 0 0 $X=188045 $Y=54965
X665 29 VIA2_C_CDNS_7246548160563 $T=188965 73955 0 0 $X=188045 $Y=73765
X666 29 VIA2_C_CDNS_7246548160563 $T=188965 92755 0 0 $X=188045 $Y=92565
X667 29 VIA2_C_CDNS_7246548160563 $T=188965 111555 0 0 $X=188045 $Y=111365
X668 29 VIA2_C_CDNS_7246548160563 $T=188965 130355 0 0 $X=188045 $Y=130165
X669 29 VIA2_C_CDNS_7246548160563 $T=188965 149155 0 0 $X=188045 $Y=148965
X670 29 VIA2_C_CDNS_7246548160563 $T=188965 167955 0 0 $X=188045 $Y=167765
X671 31 VIA2_C_CDNS_7246548160563 $T=191245 55935 0 0 $X=190325 $Y=55745
X672 31 VIA2_C_CDNS_7246548160563 $T=191245 74735 0 0 $X=190325 $Y=74545
X673 31 VIA2_C_CDNS_7246548160563 $T=191245 93535 0 0 $X=190325 $Y=93345
X674 31 VIA2_C_CDNS_7246548160563 $T=191245 112335 0 0 $X=190325 $Y=112145
X675 31 VIA2_C_CDNS_7246548160563 $T=191245 131135 0 0 $X=190325 $Y=130945
X676 31 VIA2_C_CDNS_7246548160563 $T=191245 149935 0 0 $X=190325 $Y=149745
X677 31 VIA2_C_CDNS_7246548160563 $T=191245 168735 0 0 $X=190325 $Y=168545
X678 28 VIA2_C_CDNS_7246548160563 $T=193525 56715 0 0 $X=192605 $Y=56525
X679 28 VIA2_C_CDNS_7246548160563 $T=193525 75515 0 0 $X=192605 $Y=75325
X680 28 VIA2_C_CDNS_7246548160563 $T=193525 94315 0 0 $X=192605 $Y=94125
X681 28 VIA2_C_CDNS_7246548160563 $T=193525 113115 0 0 $X=192605 $Y=112925
X682 28 VIA2_C_CDNS_7246548160563 $T=193525 131915 0 0 $X=192605 $Y=131725
X683 28 VIA2_C_CDNS_7246548160563 $T=193525 150715 0 0 $X=192605 $Y=150525
X684 28 VIA2_C_CDNS_7246548160563 $T=193525 169515 0 0 $X=192605 $Y=169325
X685 27 VIA2_C_CDNS_7246548160563 $T=195805 57495 0 0 $X=194885 $Y=57305
X686 27 VIA2_C_CDNS_7246548160563 $T=195805 76295 0 0 $X=194885 $Y=76105
X687 27 VIA2_C_CDNS_7246548160563 $T=195805 95095 0 0 $X=194885 $Y=94905
X688 27 VIA2_C_CDNS_7246548160563 $T=195805 113895 0 0 $X=194885 $Y=113705
X689 27 VIA2_C_CDNS_7246548160563 $T=195805 132695 0 0 $X=194885 $Y=132505
X690 27 VIA2_C_CDNS_7246548160563 $T=195805 151495 0 0 $X=194885 $Y=151305
X691 27 VIA2_C_CDNS_7246548160563 $T=195805 170295 0 0 $X=194885 $Y=170105
X692 26 VIA2_C_CDNS_7246548160563 $T=198085 58275 0 0 $X=197165 $Y=58085
X693 26 VIA2_C_CDNS_7246548160563 $T=198085 77075 0 0 $X=197165 $Y=76885
X694 26 VIA2_C_CDNS_7246548160563 $T=198085 95875 0 0 $X=197165 $Y=95685
X695 26 VIA2_C_CDNS_7246548160563 $T=198085 114675 0 0 $X=197165 $Y=114485
X696 26 VIA2_C_CDNS_7246548160563 $T=198085 133475 0 0 $X=197165 $Y=133285
X697 26 VIA2_C_CDNS_7246548160563 $T=198085 152275 0 0 $X=197165 $Y=152085
X698 26 VIA2_C_CDNS_7246548160563 $T=198085 171075 0 0 $X=197165 $Y=170885
X699 30 VIA2_C_CDNS_7246548160563 $T=200365 59055 0 0 $X=199445 $Y=58865
X700 30 VIA2_C_CDNS_7246548160563 $T=200365 77855 0 0 $X=199445 $Y=77665
X701 30 VIA2_C_CDNS_7246548160563 $T=200365 96655 0 0 $X=199445 $Y=96465
X702 30 VIA2_C_CDNS_7246548160563 $T=200365 115455 0 0 $X=199445 $Y=115265
X703 30 VIA2_C_CDNS_7246548160563 $T=200365 134255 0 0 $X=199445 $Y=134065
X704 30 VIA2_C_CDNS_7246548160563 $T=200365 153055 0 0 $X=199445 $Y=152865
X705 30 VIA2_C_CDNS_7246548160563 $T=200365 171855 0 0 $X=199445 $Y=171665
X706 2 VIA2_C_CDNS_7246548160563 $T=202645 48755 0 0 $X=201725 $Y=48565
X707 2 VIA2_C_CDNS_7246548160563 $T=202645 59835 0 0 $X=201725 $Y=59645
X708 2 VIA2_C_CDNS_7246548160563 $T=202645 78635 0 0 $X=201725 $Y=78445
X709 2 VIA2_C_CDNS_7246548160563 $T=202645 97435 0 0 $X=201725 $Y=97245
X710 2 VIA2_C_CDNS_7246548160563 $T=202645 116235 0 0 $X=201725 $Y=116045
X711 2 VIA2_C_CDNS_7246548160563 $T=202645 135035 0 0 $X=201725 $Y=134845
X712 2 VIA2_C_CDNS_7246548160563 $T=202645 153835 0 0 $X=201725 $Y=153645
X713 2 VIA2_C_CDNS_7246548160563 $T=202645 172635 0 0 $X=201725 $Y=172445
X714 2 VIA2_C_CDNS_7246548160563 $T=202645 177475 0 0 $X=201725 $Y=177285
X715 2 VIA2_C_CDNS_7246548160563 $T=375585 48755 0 0 $X=374665 $Y=48565
X716 2 VIA2_C_CDNS_7246548160563 $T=375585 59835 0 0 $X=374665 $Y=59645
X717 2 VIA2_C_CDNS_7246548160563 $T=375585 78635 0 0 $X=374665 $Y=78445
X718 2 VIA2_C_CDNS_7246548160563 $T=375585 97435 0 0 $X=374665 $Y=97245
X719 2 VIA2_C_CDNS_7246548160563 $T=375585 116235 0 0 $X=374665 $Y=116045
X720 2 VIA2_C_CDNS_7246548160563 $T=375585 135035 0 0 $X=374665 $Y=134845
X721 2 VIA2_C_CDNS_7246548160563 $T=375585 153835 0 0 $X=374665 $Y=153645
X722 2 VIA2_C_CDNS_7246548160563 $T=375585 172635 0 0 $X=374665 $Y=172445
X723 2 VIA2_C_CDNS_7246548160563 $T=375585 177475 0 0 $X=374665 $Y=177285
X724 24 VIA2_C_CDNS_7246548160563 $T=377865 53595 0 0 $X=376945 $Y=53405
X725 24 VIA2_C_CDNS_7246548160563 $T=377865 72395 0 0 $X=376945 $Y=72205
X726 24 VIA2_C_CDNS_7246548160563 $T=377865 91195 0 0 $X=376945 $Y=91005
X727 24 VIA2_C_CDNS_7246548160563 $T=377865 109995 0 0 $X=376945 $Y=109805
X728 24 VIA2_C_CDNS_7246548160563 $T=377865 128795 0 0 $X=376945 $Y=128605
X729 24 VIA2_C_CDNS_7246548160563 $T=377865 147595 0 0 $X=376945 $Y=147405
X730 24 VIA2_C_CDNS_7246548160563 $T=377865 166395 0 0 $X=376945 $Y=166205
X731 17 VIA2_C_CDNS_7246548160563 $T=380145 54375 0 0 $X=379225 $Y=54185
X732 17 VIA2_C_CDNS_7246548160563 $T=380145 73175 0 0 $X=379225 $Y=72985
X733 17 VIA2_C_CDNS_7246548160563 $T=380145 91975 0 0 $X=379225 $Y=91785
X734 17 VIA2_C_CDNS_7246548160563 $T=380145 110775 0 0 $X=379225 $Y=110585
X735 17 VIA2_C_CDNS_7246548160563 $T=380145 129575 0 0 $X=379225 $Y=129385
X736 17 VIA2_C_CDNS_7246548160563 $T=380145 148375 0 0 $X=379225 $Y=148185
X737 17 VIA2_C_CDNS_7246548160563 $T=380145 167175 0 0 $X=379225 $Y=166985
X738 29 VIA2_C_CDNS_7246548160563 $T=382425 55155 0 0 $X=381505 $Y=54965
X739 29 VIA2_C_CDNS_7246548160563 $T=382425 73955 0 0 $X=381505 $Y=73765
X740 29 VIA2_C_CDNS_7246548160563 $T=382425 92755 0 0 $X=381505 $Y=92565
X741 29 VIA2_C_CDNS_7246548160563 $T=382425 111555 0 0 $X=381505 $Y=111365
X742 29 VIA2_C_CDNS_7246548160563 $T=382425 130355 0 0 $X=381505 $Y=130165
X743 29 VIA2_C_CDNS_7246548160563 $T=382425 149155 0 0 $X=381505 $Y=148965
X744 29 VIA2_C_CDNS_7246548160563 $T=382425 167955 0 0 $X=381505 $Y=167765
X745 31 VIA2_C_CDNS_7246548160563 $T=384705 55935 0 0 $X=383785 $Y=55745
X746 31 VIA2_C_CDNS_7246548160563 $T=384705 74735 0 0 $X=383785 $Y=74545
X747 31 VIA2_C_CDNS_7246548160563 $T=384705 93535 0 0 $X=383785 $Y=93345
X748 31 VIA2_C_CDNS_7246548160563 $T=384705 112335 0 0 $X=383785 $Y=112145
X749 31 VIA2_C_CDNS_7246548160563 $T=384705 131135 0 0 $X=383785 $Y=130945
X750 31 VIA2_C_CDNS_7246548160563 $T=384705 149935 0 0 $X=383785 $Y=149745
X751 31 VIA2_C_CDNS_7246548160563 $T=384705 168735 0 0 $X=383785 $Y=168545
X752 28 VIA2_C_CDNS_7246548160563 $T=386985 56715 0 0 $X=386065 $Y=56525
X753 28 VIA2_C_CDNS_7246548160563 $T=386985 75515 0 0 $X=386065 $Y=75325
X754 28 VIA2_C_CDNS_7246548160563 $T=386985 94315 0 0 $X=386065 $Y=94125
X755 28 VIA2_C_CDNS_7246548160563 $T=386985 113115 0 0 $X=386065 $Y=112925
X756 28 VIA2_C_CDNS_7246548160563 $T=386985 131915 0 0 $X=386065 $Y=131725
X757 28 VIA2_C_CDNS_7246548160563 $T=386985 150715 0 0 $X=386065 $Y=150525
X758 28 VIA2_C_CDNS_7246548160563 $T=386985 169515 0 0 $X=386065 $Y=169325
X759 27 VIA2_C_CDNS_7246548160563 $T=389265 57495 0 0 $X=388345 $Y=57305
X760 27 VIA2_C_CDNS_7246548160563 $T=389265 76295 0 0 $X=388345 $Y=76105
X761 27 VIA2_C_CDNS_7246548160563 $T=389265 95095 0 0 $X=388345 $Y=94905
X762 27 VIA2_C_CDNS_7246548160563 $T=389265 113895 0 0 $X=388345 $Y=113705
X763 27 VIA2_C_CDNS_7246548160563 $T=389265 132695 0 0 $X=388345 $Y=132505
X764 27 VIA2_C_CDNS_7246548160563 $T=389265 151495 0 0 $X=388345 $Y=151305
X765 27 VIA2_C_CDNS_7246548160563 $T=389265 170295 0 0 $X=388345 $Y=170105
X766 26 VIA2_C_CDNS_7246548160563 $T=391545 58275 0 0 $X=390625 $Y=58085
X767 26 VIA2_C_CDNS_7246548160563 $T=391545 77075 0 0 $X=390625 $Y=76885
X768 26 VIA2_C_CDNS_7246548160563 $T=391545 95875 0 0 $X=390625 $Y=95685
X769 26 VIA2_C_CDNS_7246548160563 $T=391545 114675 0 0 $X=390625 $Y=114485
X770 26 VIA2_C_CDNS_7246548160563 $T=391545 133475 0 0 $X=390625 $Y=133285
X771 26 VIA2_C_CDNS_7246548160563 $T=391545 152275 0 0 $X=390625 $Y=152085
X772 26 VIA2_C_CDNS_7246548160563 $T=391545 171075 0 0 $X=390625 $Y=170885
X773 30 VIA2_C_CDNS_7246548160563 $T=393825 59055 0 0 $X=392905 $Y=58865
X774 30 VIA2_C_CDNS_7246548160563 $T=393825 77855 0 0 $X=392905 $Y=77665
X775 30 VIA2_C_CDNS_7246548160563 $T=393825 96655 0 0 $X=392905 $Y=96465
X776 30 VIA2_C_CDNS_7246548160563 $T=393825 115455 0 0 $X=392905 $Y=115265
X777 30 VIA2_C_CDNS_7246548160563 $T=393825 134255 0 0 $X=392905 $Y=134065
X778 30 VIA2_C_CDNS_7246548160563 $T=393825 153055 0 0 $X=392905 $Y=152865
X779 30 VIA2_C_CDNS_7246548160563 $T=393825 171855 0 0 $X=392905 $Y=171665
X780 30 VIA1_C_CDNS_7246548160564 $T=223665 38490 1 0 $X=223265 $Y=37520
X781 23 VIA1_C_CDNS_7246548160564 $T=225205 40770 1 0 $X=224805 $Y=39800
X782 30 VIA1_C_CDNS_7246548160564 $T=226745 38490 1 0 $X=226345 $Y=37520
X783 23 VIA1_C_CDNS_7246548160564 $T=228285 40770 1 0 $X=227885 $Y=39800
X784 30 VIA1_C_CDNS_7246548160564 $T=229825 38490 1 0 $X=229425 $Y=37520
X785 23 VIA1_C_CDNS_7246548160564 $T=231365 40770 1 0 $X=230965 $Y=39800
X786 30 VIA1_C_CDNS_7246548160564 $T=232905 38490 1 0 $X=232505 $Y=37520
X787 23 VIA1_C_CDNS_7246548160564 $T=234445 40770 1 0 $X=234045 $Y=39800
X788 30 VIA1_C_CDNS_7246548160564 $T=235985 38490 1 0 $X=235585 $Y=37520
X789 23 VIA1_C_CDNS_7246548160564 $T=237525 40770 1 0 $X=237125 $Y=39800
X790 30 VIA1_C_CDNS_7246548160564 $T=239065 38490 1 0 $X=238665 $Y=37520
X791 26 VIA1_C_CDNS_7246548160564 $T=246485 40770 1 0 $X=246085 $Y=39800
X792 5 VIA1_C_CDNS_7246548160564 $T=248025 38490 1 0 $X=247625 $Y=37520
X793 26 VIA1_C_CDNS_7246548160564 $T=249565 40770 1 0 $X=249165 $Y=39800
X794 5 VIA1_C_CDNS_7246548160564 $T=251105 38490 1 0 $X=250705 $Y=37520
X795 26 VIA1_C_CDNS_7246548160564 $T=252645 40770 1 0 $X=252245 $Y=39800
X796 5 VIA1_C_CDNS_7246548160564 $T=254185 38490 1 0 $X=253785 $Y=37520
X797 26 VIA1_C_CDNS_7246548160564 $T=255725 40770 1 0 $X=255325 $Y=39800
X798 5 VIA1_C_CDNS_7246548160564 $T=257265 38490 1 0 $X=256865 $Y=37520
X799 26 VIA1_C_CDNS_7246548160564 $T=258805 40770 1 0 $X=258405 $Y=39800
X800 5 VIA1_C_CDNS_7246548160564 $T=260345 38490 1 0 $X=259945 $Y=37520
X801 26 VIA1_C_CDNS_7246548160564 $T=261885 40770 1 0 $X=261485 $Y=39800
X802 5 VIA1_C_CDNS_7246548160564 $T=263425 38490 1 0 $X=263025 $Y=37520
X803 26 VIA1_C_CDNS_7246548160564 $T=264965 40770 1 0 $X=264565 $Y=39800
X804 5 VIA1_C_CDNS_7246548160564 $T=266505 38490 1 0 $X=266105 $Y=37520
X805 26 VIA1_C_CDNS_7246548160564 $T=268045 40770 1 0 $X=267645 $Y=39800
X806 5 VIA1_C_CDNS_7246548160564 $T=269585 38490 1 0 $X=269185 $Y=37520
X807 26 VIA1_C_CDNS_7246548160564 $T=271125 40770 1 0 $X=270725 $Y=39800
X808 5 VIA1_C_CDNS_7246548160564 $T=272665 38490 1 0 $X=272265 $Y=37520
X809 26 VIA1_C_CDNS_7246548160564 $T=274205 40770 1 0 $X=273805 $Y=39800
X810 5 VIA1_C_CDNS_7246548160564 $T=275745 38490 1 0 $X=275345 $Y=37520
X811 26 VIA1_C_CDNS_7246548160564 $T=277285 40770 1 0 $X=276885 $Y=39800
X812 5 VIA1_C_CDNS_7246548160564 $T=278825 38490 1 0 $X=278425 $Y=37520
X813 26 VIA1_C_CDNS_7246548160564 $T=280365 40770 1 0 $X=279965 $Y=39800
X814 5 VIA1_C_CDNS_7246548160564 $T=281905 38490 1 0 $X=281505 $Y=37520
X815 26 VIA1_C_CDNS_7246548160564 $T=283445 40770 1 0 $X=283045 $Y=39800
X816 5 VIA1_C_CDNS_7246548160564 $T=284985 38490 1 0 $X=284585 $Y=37520
X817 26 VIA1_C_CDNS_7246548160564 $T=286525 40770 1 0 $X=286125 $Y=39800
X818 5 VIA1_C_CDNS_7246548160564 $T=288065 38490 1 0 $X=287665 $Y=37520
X819 26 VIA1_C_CDNS_7246548160564 $T=289605 40770 1 0 $X=289205 $Y=39800
X820 5 VIA1_C_CDNS_7246548160564 $T=291145 38490 1 0 $X=290745 $Y=37520
X821 26 VIA1_C_CDNS_7246548160564 $T=292685 40770 1 0 $X=292285 $Y=39800
X822 5 VIA1_C_CDNS_7246548160564 $T=294225 38490 1 0 $X=293825 $Y=37520
X823 26 VIA1_C_CDNS_7246548160564 $T=295765 40770 1 0 $X=295365 $Y=39800
X824 27 VIA1_C_CDNS_7246548160564 $T=302300 40770 1 0 $X=301900 $Y=39800
X825 5 VIA1_C_CDNS_7246548160564 $T=303840 38490 1 0 $X=303440 $Y=37520
X826 27 VIA1_C_CDNS_7246548160564 $T=305380 40770 1 0 $X=304980 $Y=39800
X827 5 VIA1_C_CDNS_7246548160564 $T=306920 38490 1 0 $X=306520 $Y=37520
X828 27 VIA1_C_CDNS_7246548160564 $T=308460 40770 1 0 $X=308060 $Y=39800
X829 5 VIA1_C_CDNS_7246548160564 $T=310000 38490 1 0 $X=309600 $Y=37520
X830 27 VIA1_C_CDNS_7246548160564 $T=311540 40770 1 0 $X=311140 $Y=39800
X831 5 VIA1_C_CDNS_7246548160564 $T=313080 38490 1 0 $X=312680 $Y=37520
X832 27 VIA1_C_CDNS_7246548160564 $T=314620 40770 1 0 $X=314220 $Y=39800
X833 5 VIA1_C_CDNS_7246548160564 $T=316160 38490 1 0 $X=315760 $Y=37520
X834 27 VIA1_C_CDNS_7246548160564 $T=317700 40770 1 0 $X=317300 $Y=39800
X835 5 VIA1_C_CDNS_7246548160564 $T=319240 38490 1 0 $X=318840 $Y=37520
X836 27 VIA1_C_CDNS_7246548160564 $T=320780 40770 1 0 $X=320380 $Y=39800
X837 5 VIA1_C_CDNS_7246548160564 $T=322320 38490 1 0 $X=321920 $Y=37520
X838 27 VIA1_C_CDNS_7246548160564 $T=323860 40770 1 0 $X=323460 $Y=39800
X839 5 VIA1_C_CDNS_7246548160564 $T=325400 38490 1 0 $X=325000 $Y=37520
X840 27 VIA1_C_CDNS_7246548160564 $T=326940 40770 1 0 $X=326540 $Y=39800
X841 28 VIA1_C_CDNS_7246548160564 $T=333065 40770 1 0 $X=332665 $Y=39800
X842 5 VIA1_C_CDNS_7246548160564 $T=334605 38490 1 0 $X=334205 $Y=37520
X843 28 VIA1_C_CDNS_7246548160564 $T=336145 40770 1 0 $X=335745 $Y=39800
X844 5 VIA1_C_CDNS_7246548160564 $T=337685 38490 1 0 $X=337285 $Y=37520
X845 28 VIA1_C_CDNS_7246548160564 $T=339225 40770 1 0 $X=338825 $Y=39800
X846 5 VIA1_C_CDNS_7246548160564 $T=340765 38490 1 0 $X=340365 $Y=37520
X847 28 VIA1_C_CDNS_7246548160564 $T=342305 40770 1 0 $X=341905 $Y=39800
X848 5 VIA1_C_CDNS_7246548160564 $T=343845 38490 1 0 $X=343445 $Y=37520
X849 28 VIA1_C_CDNS_7246548160564 $T=345385 40770 1 0 $X=344985 $Y=39800
X850 31 VIA1_C_CDNS_7246548160564 $T=351530 40770 1 0 $X=351130 $Y=39800
X851 5 VIA1_C_CDNS_7246548160564 $T=353070 38490 1 0 $X=352670 $Y=37520
X852 31 VIA1_C_CDNS_7246548160564 $T=354610 40770 1 0 $X=354210 $Y=39800
X853 5 VIA1_C_CDNS_7246548160564 $T=356150 38490 1 0 $X=355750 $Y=37520
X854 31 VIA1_C_CDNS_7246548160564 $T=357690 40770 1 0 $X=357290 $Y=39800
X855 29 VIA1_C_CDNS_7246548160564 $T=363865 40770 1 0 $X=363465 $Y=39800
X856 5 VIA1_C_CDNS_7246548160564 $T=365405 38490 1 0 $X=365005 $Y=37520
X857 29 VIA1_C_CDNS_7246548160564 $T=366945 40770 1 0 $X=366545 $Y=39800
X858 24 VIA1_C_CDNS_7246548160564 $T=373240 40770 1 0 $X=372840 $Y=39800
X859 5 VIA1_C_CDNS_7246548160564 $T=374780 38490 1 0 $X=374380 $Y=37520
X860 15 VIA2_C_CDNS_7246548160565 $T=10890 144880 0 0 $X=10180 $Y=144220
X861 15 VIA2_C_CDNS_7246548160565 $T=10890 177040 0 0 $X=10180 $Y=176380
X862 20 VIA2_C_CDNS_7246548160565 $T=41770 143100 0 0 $X=41060 $Y=142440
X863 20 VIA2_C_CDNS_7246548160565 $T=41770 175260 0 0 $X=41060 $Y=174600
X864 2 VIA1_C_CDNS_7246548160567 $T=79820 146660 0 0 $X=78380 $Y=146470
X865 2 VIA1_C_CDNS_7246548160567 $T=79820 173480 0 0 $X=78380 $Y=173290
X866 2 VIA1_C_CDNS_7246548160567 $T=91060 146660 0 0 $X=89620 $Y=146470
X867 2 VIA1_C_CDNS_7246548160567 $T=91060 173480 0 0 $X=89620 $Y=173290
X868 2 VIA1_C_CDNS_7246548160567 $T=102300 146660 0 0 $X=100860 $Y=146470
X869 2 VIA1_C_CDNS_7246548160567 $T=102300 173480 0 0 $X=100860 $Y=173290
X870 2 VIA1_C_CDNS_7246548160567 $T=113540 146660 0 0 $X=112100 $Y=146470
X871 2 VIA1_C_CDNS_7246548160567 $T=113540 173480 0 0 $X=112100 $Y=173290
X872 2 VIA1_C_CDNS_7246548160567 $T=124780 146660 0 0 $X=123340 $Y=146470
X873 2 VIA1_C_CDNS_7246548160567 $T=124780 173480 0 0 $X=123340 $Y=173290
X874 2 VIA1_C_CDNS_7246548160567 $T=136020 146660 0 0 $X=134580 $Y=146470
X875 2 VIA1_C_CDNS_7246548160567 $T=136020 173480 0 0 $X=134580 $Y=173290
X876 2 VIA1_C_CDNS_7246548160567 $T=147260 146660 0 0 $X=145820 $Y=146470
X877 2 VIA1_C_CDNS_7246548160567 $T=147260 173480 0 0 $X=145820 $Y=173290
X878 2 VIA1_C_CDNS_7246548160567 $T=158500 146660 0 0 $X=157060 $Y=146470
X879 2 VIA1_C_CDNS_7246548160567 $T=158500 173480 0 0 $X=157060 $Y=173290
X880 22 VIA2_C_CDNS_7246548160568 $T=70100 98685 0 0 $X=69960 $Y=97975
X881 22 VIA2_C_CDNS_7246548160568 $T=70100 126585 0 0 $X=69960 $Y=125875
X882 22 VIA2_C_CDNS_7246548160568 $T=71370 98685 0 0 $X=71230 $Y=97975
X883 22 VIA2_C_CDNS_7246548160568 $T=71370 126585 0 0 $X=71230 $Y=125875
X884 22 VIA2_C_CDNS_7246548160568 $T=72640 98685 0 0 $X=72500 $Y=97975
X885 22 VIA2_C_CDNS_7246548160568 $T=72640 126585 0 0 $X=72500 $Y=125875
X886 22 VIA2_C_CDNS_7246548160568 $T=73500 98685 0 0 $X=73360 $Y=97975
X887 22 VIA2_C_CDNS_7246548160568 $T=73500 126585 0 0 $X=73360 $Y=125875
X888 22 VIA2_C_CDNS_7246548160568 $T=74770 98685 0 0 $X=74630 $Y=97975
X889 22 VIA2_C_CDNS_7246548160568 $T=74770 126585 0 0 $X=74630 $Y=125875
X890 16 VIA2_C_CDNS_7246548160568 $T=76040 96905 0 0 $X=75900 $Y=96195
X891 17 VIA2_C_CDNS_7246548160568 $T=76040 128365 0 0 $X=75900 $Y=127655
X892 22 VIA2_C_CDNS_7246548160568 $T=76900 98685 0 0 $X=76760 $Y=97975
X893 22 VIA2_C_CDNS_7246548160568 $T=76900 126585 0 0 $X=76760 $Y=125875
X894 22 VIA2_C_CDNS_7246548160568 $T=78170 98685 0 0 $X=78030 $Y=97975
X895 22 VIA2_C_CDNS_7246548160568 $T=78170 126585 0 0 $X=78030 $Y=125875
X896 17 VIA2_C_CDNS_7246548160568 $T=79440 95125 0 0 $X=79300 $Y=94415
X897 16 VIA2_C_CDNS_7246548160568 $T=79440 130145 0 0 $X=79300 $Y=129435
X898 22 VIA2_C_CDNS_7246548160568 $T=80300 98685 0 0 $X=80160 $Y=97975
X899 22 VIA2_C_CDNS_7246548160568 $T=80300 126585 0 0 $X=80160 $Y=125875
X900 22 VIA2_C_CDNS_7246548160568 $T=81570 98685 0 0 $X=81430 $Y=97975
X901 22 VIA2_C_CDNS_7246548160568 $T=81570 126585 0 0 $X=81430 $Y=125875
X902 16 VIA2_C_CDNS_7246548160568 $T=82840 96905 0 0 $X=82700 $Y=96195
X903 17 VIA2_C_CDNS_7246548160568 $T=82840 128365 0 0 $X=82700 $Y=127655
X904 22 VIA2_C_CDNS_7246548160568 $T=83700 98685 0 0 $X=83560 $Y=97975
X905 22 VIA2_C_CDNS_7246548160568 $T=83700 126585 0 0 $X=83560 $Y=125875
X906 22 VIA2_C_CDNS_7246548160568 $T=84970 98685 0 0 $X=84830 $Y=97975
X907 22 VIA2_C_CDNS_7246548160568 $T=84970 126585 0 0 $X=84830 $Y=125875
X908 17 VIA2_C_CDNS_7246548160568 $T=86240 95125 0 0 $X=86100 $Y=94415
X909 16 VIA2_C_CDNS_7246548160568 $T=86240 130145 0 0 $X=86100 $Y=129435
X910 22 VIA2_C_CDNS_7246548160568 $T=87100 98685 0 0 $X=86960 $Y=97975
X911 22 VIA2_C_CDNS_7246548160568 $T=87100 126585 0 0 $X=86960 $Y=125875
X912 22 VIA2_C_CDNS_7246548160568 $T=88370 98685 0 0 $X=88230 $Y=97975
X913 22 VIA2_C_CDNS_7246548160568 $T=88370 126585 0 0 $X=88230 $Y=125875
X914 16 VIA2_C_CDNS_7246548160568 $T=89640 96905 0 0 $X=89500 $Y=96195
X915 17 VIA2_C_CDNS_7246548160568 $T=89640 128365 0 0 $X=89500 $Y=127655
X916 22 VIA2_C_CDNS_7246548160568 $T=90500 98685 0 0 $X=90360 $Y=97975
X917 22 VIA2_C_CDNS_7246548160568 $T=90500 126585 0 0 $X=90360 $Y=125875
X918 22 VIA2_C_CDNS_7246548160568 $T=91770 98685 0 0 $X=91630 $Y=97975
X919 22 VIA2_C_CDNS_7246548160568 $T=91770 126585 0 0 $X=91630 $Y=125875
X920 17 VIA2_C_CDNS_7246548160568 $T=93040 95125 0 0 $X=92900 $Y=94415
X921 16 VIA2_C_CDNS_7246548160568 $T=93040 130145 0 0 $X=92900 $Y=129435
X922 22 VIA2_C_CDNS_7246548160568 $T=93900 98685 0 0 $X=93760 $Y=97975
X923 22 VIA2_C_CDNS_7246548160568 $T=93900 126585 0 0 $X=93760 $Y=125875
X924 22 VIA2_C_CDNS_7246548160568 $T=95170 98685 0 0 $X=95030 $Y=97975
X925 22 VIA2_C_CDNS_7246548160568 $T=95170 126585 0 0 $X=95030 $Y=125875
X926 16 VIA2_C_CDNS_7246548160568 $T=96440 96905 0 0 $X=96300 $Y=96195
X927 17 VIA2_C_CDNS_7246548160568 $T=96440 128365 0 0 $X=96300 $Y=127655
X928 22 VIA2_C_CDNS_7246548160568 $T=97300 98685 0 0 $X=97160 $Y=97975
X929 22 VIA2_C_CDNS_7246548160568 $T=97300 126585 0 0 $X=97160 $Y=125875
X930 22 VIA2_C_CDNS_7246548160568 $T=98570 98685 0 0 $X=98430 $Y=97975
X931 22 VIA2_C_CDNS_7246548160568 $T=98570 126585 0 0 $X=98430 $Y=125875
X932 17 VIA2_C_CDNS_7246548160568 $T=99840 95125 0 0 $X=99700 $Y=94415
X933 16 VIA2_C_CDNS_7246548160568 $T=99840 130145 0 0 $X=99700 $Y=129435
X934 22 VIA2_C_CDNS_7246548160568 $T=100700 98685 0 0 $X=100560 $Y=97975
X935 22 VIA2_C_CDNS_7246548160568 $T=100700 126585 0 0 $X=100560 $Y=125875
X936 22 VIA2_C_CDNS_7246548160568 $T=101970 98685 0 0 $X=101830 $Y=97975
X937 22 VIA2_C_CDNS_7246548160568 $T=101970 126585 0 0 $X=101830 $Y=125875
X938 16 VIA2_C_CDNS_7246548160568 $T=103240 96905 0 0 $X=103100 $Y=96195
X939 17 VIA2_C_CDNS_7246548160568 $T=103240 128365 0 0 $X=103100 $Y=127655
X940 22 VIA2_C_CDNS_7246548160568 $T=104100 98685 0 0 $X=103960 $Y=97975
X941 22 VIA2_C_CDNS_7246548160568 $T=104100 126585 0 0 $X=103960 $Y=125875
X942 22 VIA2_C_CDNS_7246548160568 $T=105370 98685 0 0 $X=105230 $Y=97975
X943 22 VIA2_C_CDNS_7246548160568 $T=105370 126585 0 0 $X=105230 $Y=125875
X944 17 VIA2_C_CDNS_7246548160568 $T=106640 95125 0 0 $X=106500 $Y=94415
X945 16 VIA2_C_CDNS_7246548160568 $T=106640 130145 0 0 $X=106500 $Y=129435
X946 22 VIA2_C_CDNS_7246548160568 $T=107500 98685 0 0 $X=107360 $Y=97975
X947 22 VIA2_C_CDNS_7246548160568 $T=107500 126585 0 0 $X=107360 $Y=125875
X948 22 VIA2_C_CDNS_7246548160568 $T=108770 98685 0 0 $X=108630 $Y=97975
X949 22 VIA2_C_CDNS_7246548160568 $T=108770 126585 0 0 $X=108630 $Y=125875
X950 16 VIA2_C_CDNS_7246548160568 $T=110040 96905 0 0 $X=109900 $Y=96195
X951 17 VIA2_C_CDNS_7246548160568 $T=110040 128365 0 0 $X=109900 $Y=127655
X952 22 VIA2_C_CDNS_7246548160568 $T=110900 98685 0 0 $X=110760 $Y=97975
X953 22 VIA2_C_CDNS_7246548160568 $T=110900 126585 0 0 $X=110760 $Y=125875
X954 22 VIA2_C_CDNS_7246548160568 $T=112170 98685 0 0 $X=112030 $Y=97975
X955 22 VIA2_C_CDNS_7246548160568 $T=112170 126585 0 0 $X=112030 $Y=125875
X956 17 VIA2_C_CDNS_7246548160568 $T=113440 95125 0 0 $X=113300 $Y=94415
X957 16 VIA2_C_CDNS_7246548160568 $T=113440 130145 0 0 $X=113300 $Y=129435
X958 22 VIA2_C_CDNS_7246548160568 $T=114300 98685 0 0 $X=114160 $Y=97975
X959 22 VIA2_C_CDNS_7246548160568 $T=114300 126585 0 0 $X=114160 $Y=125875
X960 22 VIA2_C_CDNS_7246548160568 $T=115570 98685 0 0 $X=115430 $Y=97975
X961 22 VIA2_C_CDNS_7246548160568 $T=115570 126585 0 0 $X=115430 $Y=125875
X962 16 VIA2_C_CDNS_7246548160568 $T=116840 96905 0 0 $X=116700 $Y=96195
X963 17 VIA2_C_CDNS_7246548160568 $T=116840 128365 0 0 $X=116700 $Y=127655
X964 22 VIA2_C_CDNS_7246548160568 $T=117700 98685 0 0 $X=117560 $Y=97975
X965 22 VIA2_C_CDNS_7246548160568 $T=117700 126585 0 0 $X=117560 $Y=125875
X966 22 VIA2_C_CDNS_7246548160568 $T=118970 98685 0 0 $X=118830 $Y=97975
X967 22 VIA2_C_CDNS_7246548160568 $T=118970 126585 0 0 $X=118830 $Y=125875
X968 17 VIA2_C_CDNS_7246548160568 $T=120240 95125 0 0 $X=120100 $Y=94415
X969 16 VIA2_C_CDNS_7246548160568 $T=120240 130145 0 0 $X=120100 $Y=129435
X970 22 VIA2_C_CDNS_7246548160568 $T=121100 98685 0 0 $X=120960 $Y=97975
X971 22 VIA2_C_CDNS_7246548160568 $T=121100 126585 0 0 $X=120960 $Y=125875
X972 22 VIA2_C_CDNS_7246548160568 $T=122370 98685 0 0 $X=122230 $Y=97975
X973 22 VIA2_C_CDNS_7246548160568 $T=122370 126585 0 0 $X=122230 $Y=125875
X974 16 VIA2_C_CDNS_7246548160568 $T=123640 96905 0 0 $X=123500 $Y=96195
X975 17 VIA2_C_CDNS_7246548160568 $T=123640 128365 0 0 $X=123500 $Y=127655
X976 22 VIA2_C_CDNS_7246548160568 $T=124500 98685 0 0 $X=124360 $Y=97975
X977 22 VIA2_C_CDNS_7246548160568 $T=124500 126585 0 0 $X=124360 $Y=125875
X978 22 VIA2_C_CDNS_7246548160568 $T=125770 98685 0 0 $X=125630 $Y=97975
X979 22 VIA2_C_CDNS_7246548160568 $T=125770 126585 0 0 $X=125630 $Y=125875
X980 17 VIA2_C_CDNS_7246548160568 $T=127040 95125 0 0 $X=126900 $Y=94415
X981 16 VIA2_C_CDNS_7246548160568 $T=127040 130145 0 0 $X=126900 $Y=129435
X982 22 VIA2_C_CDNS_7246548160568 $T=127900 98685 0 0 $X=127760 $Y=97975
X983 22 VIA2_C_CDNS_7246548160568 $T=127900 126585 0 0 $X=127760 $Y=125875
X984 22 VIA2_C_CDNS_7246548160568 $T=129170 98685 0 0 $X=129030 $Y=97975
X985 22 VIA2_C_CDNS_7246548160568 $T=129170 126585 0 0 $X=129030 $Y=125875
X986 22 VIA2_C_CDNS_7246548160568 $T=130440 98685 0 0 $X=130300 $Y=97975
X987 22 VIA2_C_CDNS_7246548160568 $T=130440 126585 0 0 $X=130300 $Y=125875
X988 22 VIA1_C_CDNS_7246548160569 $T=71370 100245 0 0 $X=70920 $Y=100105
X989 22 VIA1_C_CDNS_7246548160569 $T=71370 125025 0 0 $X=70920 $Y=124885
X990 22 VIA1_C_CDNS_7246548160569 $T=74770 100245 0 0 $X=74320 $Y=100105
X991 22 VIA1_C_CDNS_7246548160569 $T=74770 125025 0 0 $X=74320 $Y=124885
X992 22 VIA1_C_CDNS_7246548160569 $T=78170 100245 0 0 $X=77720 $Y=100105
X993 22 VIA1_C_CDNS_7246548160569 $T=78170 125025 0 0 $X=77720 $Y=124885
X994 22 VIA1_C_CDNS_7246548160569 $T=81570 100245 0 0 $X=81120 $Y=100105
X995 22 VIA1_C_CDNS_7246548160569 $T=81570 125025 0 0 $X=81120 $Y=124885
X996 22 VIA1_C_CDNS_7246548160569 $T=84970 100245 0 0 $X=84520 $Y=100105
X997 22 VIA1_C_CDNS_7246548160569 $T=84970 125025 0 0 $X=84520 $Y=124885
X998 22 VIA1_C_CDNS_7246548160569 $T=88370 100245 0 0 $X=87920 $Y=100105
X999 22 VIA1_C_CDNS_7246548160569 $T=88370 125025 0 0 $X=87920 $Y=124885
X1000 22 VIA1_C_CDNS_7246548160569 $T=91770 100245 0 0 $X=91320 $Y=100105
X1001 22 VIA1_C_CDNS_7246548160569 $T=91770 125025 0 0 $X=91320 $Y=124885
X1002 22 VIA1_C_CDNS_7246548160569 $T=95170 100245 0 0 $X=94720 $Y=100105
X1003 22 VIA1_C_CDNS_7246548160569 $T=95170 125025 0 0 $X=94720 $Y=124885
X1004 22 VIA1_C_CDNS_7246548160569 $T=98570 100245 0 0 $X=98120 $Y=100105
X1005 22 VIA1_C_CDNS_7246548160569 $T=98570 125025 0 0 $X=98120 $Y=124885
X1006 22 VIA1_C_CDNS_7246548160569 $T=101970 100245 0 0 $X=101520 $Y=100105
X1007 22 VIA1_C_CDNS_7246548160569 $T=101970 125025 0 0 $X=101520 $Y=124885
X1008 22 VIA1_C_CDNS_7246548160569 $T=105370 100245 0 0 $X=104920 $Y=100105
X1009 22 VIA1_C_CDNS_7246548160569 $T=105370 125025 0 0 $X=104920 $Y=124885
X1010 22 VIA1_C_CDNS_7246548160569 $T=108770 100245 0 0 $X=108320 $Y=100105
X1011 22 VIA1_C_CDNS_7246548160569 $T=108770 125025 0 0 $X=108320 $Y=124885
X1012 22 VIA1_C_CDNS_7246548160569 $T=112170 100245 0 0 $X=111720 $Y=100105
X1013 22 VIA1_C_CDNS_7246548160569 $T=112170 125025 0 0 $X=111720 $Y=124885
X1014 22 VIA1_C_CDNS_7246548160569 $T=115570 100245 0 0 $X=115120 $Y=100105
X1015 22 VIA1_C_CDNS_7246548160569 $T=115570 125025 0 0 $X=115120 $Y=124885
X1016 22 VIA1_C_CDNS_7246548160569 $T=118970 100245 0 0 $X=118520 $Y=100105
X1017 22 VIA1_C_CDNS_7246548160569 $T=118970 125025 0 0 $X=118520 $Y=124885
X1018 22 VIA1_C_CDNS_7246548160569 $T=122370 100245 0 0 $X=121920 $Y=100105
X1019 22 VIA1_C_CDNS_7246548160569 $T=122370 125025 0 0 $X=121920 $Y=124885
X1020 22 VIA1_C_CDNS_7246548160569 $T=125770 100245 0 0 $X=125320 $Y=100105
X1021 22 VIA1_C_CDNS_7246548160569 $T=125770 125025 0 0 $X=125320 $Y=124885
X1022 22 VIA1_C_CDNS_7246548160569 $T=129170 100245 0 0 $X=128720 $Y=100105
X1023 22 VIA1_C_CDNS_7246548160569 $T=129170 125025 0 0 $X=128720 $Y=124885
X1024 17 VIA3_C_CDNS_7246548160570 $T=63650 95125 0 0 $X=62680 $Y=94465
X1025 17 VIA3_C_CDNS_7246548160570 $T=63650 128365 0 0 $X=62680 $Y=127705
X1026 16 VIA3_C_CDNS_7246548160570 $T=65930 96905 0 0 $X=64960 $Y=96245
X1027 16 VIA3_C_CDNS_7246548160570 $T=65930 130145 0 0 $X=64960 $Y=129485
X1028 22 VIA3_C_CDNS_7246548160570 $T=68210 98685 0 0 $X=67240 $Y=98025
X1029 22 VIA3_C_CDNS_7246548160570 $T=68210 126585 0 0 $X=67240 $Y=125925
X1030 22 VIA3_C_CDNS_7246548160570 $T=132330 98685 0 0 $X=131360 $Y=98025
X1031 22 VIA3_C_CDNS_7246548160570 $T=132330 126585 0 0 $X=131360 $Y=125925
X1032 17 VIA3_C_CDNS_7246548160570 $T=134610 95125 0 0 $X=133640 $Y=94465
X1033 17 VIA3_C_CDNS_7246548160570 $T=134610 128365 0 0 $X=133640 $Y=127705
X1034 16 VIA3_C_CDNS_7246548160570 $T=136890 96905 0 0 $X=135920 $Y=96245
X1035 16 VIA3_C_CDNS_7246548160570 $T=136890 130145 0 0 $X=135920 $Y=129485
X1036 6 VIA2_C_CDNS_7246548160571 $T=74460 112235 0 0 $X=74320 $Y=112045
X1037 23 VIA2_C_CDNS_7246548160571 $T=75080 113015 0 0 $X=74940 $Y=112825
X1038 6 VIA2_C_CDNS_7246548160571 $T=78170 112235 0 0 $X=78030 $Y=112045
X1039 23 VIA2_C_CDNS_7246548160571 $T=78170 113015 0 0 $X=78030 $Y=112825
X1040 6 VIA2_C_CDNS_7246548160571 $T=81260 112235 0 0 $X=81120 $Y=112045
X1041 23 VIA2_C_CDNS_7246548160571 $T=81880 113015 0 0 $X=81740 $Y=112825
X1042 6 VIA2_C_CDNS_7246548160571 $T=84970 112235 0 0 $X=84830 $Y=112045
X1043 23 VIA2_C_CDNS_7246548160571 $T=84970 113015 0 0 $X=84830 $Y=112825
X1044 6 VIA2_C_CDNS_7246548160571 $T=88060 112235 0 0 $X=87920 $Y=112045
X1045 23 VIA2_C_CDNS_7246548160571 $T=88680 113015 0 0 $X=88540 $Y=112825
X1046 6 VIA2_C_CDNS_7246548160571 $T=91770 112235 0 0 $X=91630 $Y=112045
X1047 23 VIA2_C_CDNS_7246548160571 $T=91770 113015 0 0 $X=91630 $Y=112825
X1048 6 VIA2_C_CDNS_7246548160571 $T=94860 112235 0 0 $X=94720 $Y=112045
X1049 23 VIA2_C_CDNS_7246548160571 $T=95480 113015 0 0 $X=95340 $Y=112825
X1050 6 VIA2_C_CDNS_7246548160571 $T=98570 112235 0 0 $X=98430 $Y=112045
X1051 23 VIA2_C_CDNS_7246548160571 $T=98570 113015 0 0 $X=98430 $Y=112825
X1052 6 VIA2_C_CDNS_7246548160571 $T=101660 112235 0 0 $X=101520 $Y=112045
X1053 23 VIA2_C_CDNS_7246548160571 $T=102280 113015 0 0 $X=102140 $Y=112825
X1054 6 VIA2_C_CDNS_7246548160571 $T=105370 112235 0 0 $X=105230 $Y=112045
X1055 23 VIA2_C_CDNS_7246548160571 $T=105370 113015 0 0 $X=105230 $Y=112825
X1056 6 VIA2_C_CDNS_7246548160571 $T=108460 112235 0 0 $X=108320 $Y=112045
X1057 23 VIA2_C_CDNS_7246548160571 $T=109080 113015 0 0 $X=108940 $Y=112825
X1058 6 VIA2_C_CDNS_7246548160571 $T=112170 112235 0 0 $X=112030 $Y=112045
X1059 23 VIA2_C_CDNS_7246548160571 $T=112170 113015 0 0 $X=112030 $Y=112825
X1060 6 VIA2_C_CDNS_7246548160571 $T=115260 112235 0 0 $X=115120 $Y=112045
X1061 23 VIA2_C_CDNS_7246548160571 $T=115880 113015 0 0 $X=115740 $Y=112825
X1062 6 VIA2_C_CDNS_7246548160571 $T=118970 112235 0 0 $X=118830 $Y=112045
X1063 23 VIA2_C_CDNS_7246548160571 $T=118970 113015 0 0 $X=118830 $Y=112825
X1064 6 VIA2_C_CDNS_7246548160571 $T=122060 112235 0 0 $X=121920 $Y=112045
X1065 23 VIA2_C_CDNS_7246548160571 $T=122680 113015 0 0 $X=122540 $Y=112825
X1066 6 VIA2_C_CDNS_7246548160571 $T=125770 112235 0 0 $X=125630 $Y=112045
X1067 23 VIA2_C_CDNS_7246548160571 $T=125770 113015 0 0 $X=125630 $Y=112825
X1068 1 VIA1_C_CDNS_7246548160573 $T=300690 18770 0 0 $X=299160 $Y=17760
X1069 1 VIA1_C_CDNS_7246548160573 $T=306120 19025 0 0 $X=304590 $Y=18015
X1070 3 VIA2_C_CDNS_7246548160574 $T=7140 58145 0 0 $X=5610 $Y=57395
X1071 13 VIA2_C_CDNS_7246548160574 $T=17075 56365 0 0 $X=15545 $Y=55615
X1072 2 1 VIA1_C_CDNS_7246548160575 $T=13915 179845 0 0 $X=8745 $Y=178835
X1073 2 1 VIA1_C_CDNS_7246548160575 $T=38730 179845 0 0 $X=33560 $Y=178835
X1074 2 1 VIA1_C_CDNS_7246548160575 $T=54060 179845 0 0 $X=48890 $Y=178835
X1075 2 1 VIA1_C_CDNS_7246548160575 $T=169780 179845 0 0 $X=164610 $Y=178835
X1076 2 1 VIA1_C_CDNS_7246548160575 $T=202645 179775 0 0 $X=197475 $Y=178765
X1077 2 1 VIA1_C_CDNS_7246548160575 $T=375600 179775 0 0 $X=370430 $Y=178765
X1078 2 1 VIA2_C_CDNS_7246548160576 $T=202645 179775 0 0 $X=197475 $Y=178765
X1079 2 1 VIA2_C_CDNS_7246548160576 $T=375600 179775 0 0 $X=370430 $Y=178765
X1080 2 VIA1_C_CDNS_7246548160577 $T=57370 119810 0 0 $X=56880 $Y=116720
X1081 2 VIA1_C_CDNS_7246548160577 $T=67590 119810 0 0 $X=67100 $Y=116720
X1082 2 VIA1_C_CDNS_7246548160577 $T=132950 119810 0 0 $X=132460 $Y=116720
X1083 2 VIA1_C_CDNS_7246548160577 $T=143170 119810 0 0 $X=142680 $Y=116720
X1084 30 VIA2_C_CDNS_7246548160580 $T=225125 38490 0 0 $X=224125 $Y=37490
X1085 26 VIA2_C_CDNS_7246548160580 $T=305715 12525 0 0 $X=304715 $Y=11525
X1086 27 VIA2_C_CDNS_7246548160580 $T=318935 12525 0 0 $X=317935 $Y=11525
X1087 28 VIA2_C_CDNS_7246548160580 $T=328195 12525 0 0 $X=327195 $Y=11525
X1088 31 VIA2_C_CDNS_7246548160580 $T=337455 12525 0 0 $X=336455 $Y=11525
X1089 29 VIA2_C_CDNS_7246548160580 $T=346715 12525 0 0 $X=345715 $Y=11525
X1090 24 VIA2_C_CDNS_7246548160580 $T=355975 12525 0 0 $X=354975 $Y=11525
X1091 21 VIA2_C_CDNS_7246548160581 $T=63460 55465 0 0 $X=61410 $Y=54455
X1092 5 VIA2_C_CDNS_7246548160581 $T=247295 38480 0 0 $X=245245 $Y=37470
X1093 26 VIA2_C_CDNS_7246548160581 $T=294955 40780 0 0 $X=292905 $Y=39770
X1094 27 VIA2_C_CDNS_7246548160581 $T=303110 40780 0 0 $X=301060 $Y=39770
X1095 28 VIA2_C_CDNS_7246548160581 $T=344575 40780 0 0 $X=342525 $Y=39770
X1096 31 VIA2_C_CDNS_7246548160581 $T=356880 40780 0 0 $X=354830 $Y=39770
X1097 29 VIA2_C_CDNS_7246548160581 $T=365495 40780 0 0 $X=363445 $Y=39770
X1098 24 VIA2_C_CDNS_7246548160581 $T=374005 40780 0 0 $X=371955 $Y=39770
X1099 27 VIA3_C_CDNS_7246548160584 $T=303110 40780 0 0 $X=301060 $Y=39770
X1100 28 VIA3_C_CDNS_7246548160584 $T=344575 40780 0 0 $X=342525 $Y=39770
X1101 24 VIA3_C_CDNS_7246548160584 $T=374005 40780 0 0 $X=371955 $Y=39770
X1102 27 VIA3_C_CDNS_7246548160586 $T=195805 49055 0 0 $X=194805 $Y=48055
X1103 24 VIA3_C_CDNS_7246548160586 $T=377865 50400 0 0 $X=376865 $Y=49400
X1104 28 VIA3_C_CDNS_7246548160586 $T=386985 47530 0 0 $X=385985 $Y=46530
X1105 18 VIA1_C_CDNS_7246548160588 $T=151480 80915 0 0 $X=150730 $Y=78865
X1106 20 VIA1_C_CDNS_7246548160588 $T=151480 122460 0 0 $X=150730 $Y=120410
X1107 2 15 15 1 pe3_CDNS_7246548160523 $T=15710 148580 0 0 $X=14200 $Y=147550
X1108 2 15 20 1 pe3_CDNS_7246548160523 $T=15710 171560 1 0 $X=14200 $Y=160530
X1109 2 15 20 1 pe3_CDNS_7246548160523 $T=26950 148580 0 0 $X=25440 $Y=147550
X1110 2 15 15 1 pe3_CDNS_7246548160523 $T=26950 171560 1 0 $X=25440 $Y=160530
X1111 2 2 2 1 pe3_CDNS_7246548160523 $T=56340 148580 0 0 $X=54830 $Y=147550
X1112 2 16 16 1 pe3_CDNS_7246548160523 $T=67580 148580 0 0 $X=66070 $Y=147550
X1113 2 16 17 1 pe3_CDNS_7246548160523 $T=78820 148580 0 0 $X=77310 $Y=147550
X1114 2 16 16 1 pe3_CDNS_7246548160523 $T=90060 148580 0 0 $X=88550 $Y=147550
X1115 2 16 17 1 pe3_CDNS_7246548160523 $T=101300 148580 0 0 $X=99790 $Y=147550
X1116 2 16 16 1 pe3_CDNS_7246548160523 $T=112540 148580 0 0 $X=111030 $Y=147550
X1117 2 16 17 1 pe3_CDNS_7246548160523 $T=123780 148580 0 0 $X=122270 $Y=147550
X1118 2 16 16 1 pe3_CDNS_7246548160523 $T=135020 148580 0 0 $X=133510 $Y=147550
X1119 2 16 17 1 pe3_CDNS_7246548160523 $T=146260 148580 0 0 $X=144750 $Y=147550
X1120 2 16 16 1 pe3_CDNS_7246548160523 $T=146260 171560 1 0 $X=144750 $Y=160530
X1121 2 2 2 1 pe3_CDNS_7246548160523 $T=157500 148580 0 0 $X=155990 $Y=147550
X1122 2 2 2 1 pe3_CDNS_7246548160523 $T=157500 171560 1 0 $X=155990 $Y=160530
X1123 2 2 2 1 pe3_CDNS_7246548160523 $T=340315 71115 1 0 $X=338805 $Y=60085
X1124 2 17 26 1 pe3_CDNS_7246548160523 $T=340315 89915 1 0 $X=338805 $Y=78885
X1125 2 17 26 1 pe3_CDNS_7246548160523 $T=340315 108715 1 0 $X=338805 $Y=97685
X1126 2 17 26 1 pe3_CDNS_7246548160523 $T=340315 127515 1 0 $X=338805 $Y=116485
X1127 2 17 26 1 pe3_CDNS_7246548160523 $T=340315 146315 1 0 $X=338805 $Y=135285
X1128 2 17 26 1 pe3_CDNS_7246548160523 $T=340315 165115 1 0 $X=338805 $Y=154085
X1129 2 2 2 1 pe3_CDNS_7246548160523 $T=351555 71115 1 0 $X=350045 $Y=60085
X1130 2 17 26 1 pe3_CDNS_7246548160523 $T=351555 89915 1 0 $X=350045 $Y=78885
X1131 2 17 26 1 pe3_CDNS_7246548160523 $T=351555 108715 1 0 $X=350045 $Y=97685
X1132 2 17 26 1 pe3_CDNS_7246548160523 $T=351555 127515 1 0 $X=350045 $Y=116485
X1133 2 17 26 1 pe3_CDNS_7246548160523 $T=351555 146315 1 0 $X=350045 $Y=135285
X1134 2 17 26 1 pe3_CDNS_7246548160523 $T=351555 165115 1 0 $X=350045 $Y=154085
X1135 2 2 2 1 pe3_CDNS_7246548160523 $T=362795 71115 1 0 $X=361285 $Y=60085
X1136 2 2 2 1 pe3_CDNS_7246548160523 $T=362795 89915 1 0 $X=361285 $Y=78885
X1137 2 2 2 1 pe3_CDNS_7246548160523 $T=362795 108715 1 0 $X=361285 $Y=97685
X1138 2 2 2 1 pe3_CDNS_7246548160523 $T=362795 127515 1 0 $X=361285 $Y=116485
X1139 2 2 2 1 pe3_CDNS_7246548160523 $T=362795 146315 1 0 $X=361285 $Y=135285
X1140 2 2 2 1 pe3_CDNS_7246548160523 $T=362795 165115 1 0 $X=361285 $Y=154085
X1141 29 19 5 2 1 pe3_CDNS_7246548160524 $T=364135 36320 1 0 $X=362625 $Y=25290
X1142 31 19 5 2 1 pe3_CDNS_7246548160525 $T=351800 36320 1 0 $X=350290 $Y=25290
X1143 28 19 5 2 1 pe3_CDNS_7246548160526 $T=333335 36320 1 0 $X=331825 $Y=25290
X1144 27 19 5 2 1 pe3_CDNS_7246548160527 $T=302570 36320 1 0 $X=301060 $Y=25290
X1145 26 19 5 2 1 pe3_CDNS_7246548160528 $T=246755 36320 1 0 $X=245245 $Y=25290
X1146 5 1 rpp1k1_3_CDNS_7246548160529 $T=190390 9160 0 0 $X=185230 $Y=8940
X1147 30 19 23 2 1 pe3_CDNS_7246548160530 $T=223935 36320 1 0 $X=222425 $Y=25290
X1148 23 1 rpp1k1_3_CDNS_7246548160531 $T=80195 9200 0 0 $X=75035 $Y=8980
X1149 18 1 1 pe3_CDNS_7246548160532 $T=154675 76695 0 0 $X=153165 $Y=75665
X1150 19 18 1 pe3_CDNS_7246548160532 $T=154675 98175 0 0 $X=153165 $Y=97145
X1151 20 19 1 pe3_CDNS_7246548160532 $T=154675 119125 0 0 $X=153165 $Y=118095
X1152 2 4 25 1 pe3_CDNS_7246548160533 $T=91085 67915 1 0 $X=90175 $Y=61345
X1153 26 7 1 2 pe3_CDNS_7246548160534 $T=307075 17335 1 0 $X=305565 $Y=6305
X1154 27 8 1 2 pe3_CDNS_7246548160534 $T=316335 17335 1 0 $X=314825 $Y=6305
X1155 28 9 1 2 pe3_CDNS_7246548160534 $T=325595 17335 1 0 $X=324085 $Y=6305
X1156 31 10 1 2 pe3_CDNS_7246548160534 $T=334855 17335 1 0 $X=333345 $Y=6305
X1157 29 11 1 2 pe3_CDNS_7246548160534 $T=344115 17335 1 0 $X=342605 $Y=6305
X1158 24 12 1 2 pe3_CDNS_7246548160534 $T=353375 17335 1 0 $X=351865 $Y=6305
X1159 13 3 3 1 ne3_CDNS_7246548160535 $T=7715 59435 0 0 $X=6915 $Y=59035
X1160 14 3 15 1 ne3_CDNS_7246548160535 $T=34470 59435 0 0 $X=33670 $Y=59035
X1161 21 3 22 1 ne3_CDNS_7246548160535 $T=62205 59435 0 0 $X=61405 $Y=59035
X1162 22 22 22 2 1 ne3i_6_CDNS_7246548160536 $T=70370 100985 0 0 $X=66310 $Y=96535
X1163 22 22 22 2 1 ne3i_6_CDNS_7246548160536 $T=70370 124285 1 0 $X=66310 $Y=109715
X1164 22 23 16 2 1 ne3i_6_CDNS_7246548160536 $T=73770 100985 0 0 $X=69710 $Y=96535
X1165 22 6 17 2 1 ne3i_6_CDNS_7246548160536 $T=73770 124285 1 0 $X=69710 $Y=109715
X1166 22 6 17 2 1 ne3i_6_CDNS_7246548160536 $T=77170 100985 0 0 $X=73110 $Y=96535
X1167 22 23 16 2 1 ne3i_6_CDNS_7246548160536 $T=77170 124285 1 0 $X=73110 $Y=109715
X1168 22 23 16 2 1 ne3i_6_CDNS_7246548160536 $T=80570 100985 0 0 $X=76510 $Y=96535
X1169 22 6 17 2 1 ne3i_6_CDNS_7246548160536 $T=80570 124285 1 0 $X=76510 $Y=109715
X1170 22 6 17 2 1 ne3i_6_CDNS_7246548160536 $T=83970 100985 0 0 $X=79910 $Y=96535
X1171 22 23 16 2 1 ne3i_6_CDNS_7246548160536 $T=83970 124285 1 0 $X=79910 $Y=109715
X1172 22 23 16 2 1 ne3i_6_CDNS_7246548160536 $T=87370 100985 0 0 $X=83310 $Y=96535
X1173 22 6 17 2 1 ne3i_6_CDNS_7246548160536 $T=87370 124285 1 0 $X=83310 $Y=109715
X1174 22 6 17 2 1 ne3i_6_CDNS_7246548160536 $T=90770 100985 0 0 $X=86710 $Y=96535
X1175 22 23 16 2 1 ne3i_6_CDNS_7246548160536 $T=90770 124285 1 0 $X=86710 $Y=109715
X1176 22 23 16 2 1 ne3i_6_CDNS_7246548160536 $T=94170 100985 0 0 $X=90110 $Y=96535
X1177 22 6 17 2 1 ne3i_6_CDNS_7246548160536 $T=94170 124285 1 0 $X=90110 $Y=109715
X1178 22 6 17 2 1 ne3i_6_CDNS_7246548160536 $T=97570 100985 0 0 $X=93510 $Y=96535
X1179 22 23 16 2 1 ne3i_6_CDNS_7246548160536 $T=97570 124285 1 0 $X=93510 $Y=109715
X1180 22 23 16 2 1 ne3i_6_CDNS_7246548160536 $T=100970 100985 0 0 $X=96910 $Y=96535
X1181 22 6 17 2 1 ne3i_6_CDNS_7246548160536 $T=100970 124285 1 0 $X=96910 $Y=109715
X1182 22 6 17 2 1 ne3i_6_CDNS_7246548160536 $T=104370 100985 0 0 $X=100310 $Y=96535
X1183 22 23 16 2 1 ne3i_6_CDNS_7246548160536 $T=104370 124285 1 0 $X=100310 $Y=109715
X1184 22 23 16 2 1 ne3i_6_CDNS_7246548160536 $T=107770 100985 0 0 $X=103710 $Y=96535
X1185 22 6 17 2 1 ne3i_6_CDNS_7246548160536 $T=107770 124285 1 0 $X=103710 $Y=109715
X1186 22 6 17 2 1 ne3i_6_CDNS_7246548160536 $T=111170 100985 0 0 $X=107110 $Y=96535
X1187 22 23 16 2 1 ne3i_6_CDNS_7246548160536 $T=111170 124285 1 0 $X=107110 $Y=109715
X1188 22 23 16 2 1 ne3i_6_CDNS_7246548160536 $T=114570 100985 0 0 $X=110510 $Y=96535
X1189 22 6 17 2 1 ne3i_6_CDNS_7246548160536 $T=114570 124285 1 0 $X=110510 $Y=109715
X1190 22 6 17 2 1 ne3i_6_CDNS_7246548160536 $T=117970 100985 0 0 $X=113910 $Y=96535
X1191 22 23 16 2 1 ne3i_6_CDNS_7246548160536 $T=117970 124285 1 0 $X=113910 $Y=109715
X1192 22 23 16 2 1 ne3i_6_CDNS_7246548160536 $T=121370 100985 0 0 $X=117310 $Y=96535
X1193 22 6 17 2 1 ne3i_6_CDNS_7246548160536 $T=121370 124285 1 0 $X=117310 $Y=109715
X1194 22 6 17 2 1 ne3i_6_CDNS_7246548160536 $T=124770 100985 0 0 $X=120710 $Y=96535
X1195 22 23 16 2 1 ne3i_6_CDNS_7246548160536 $T=124770 124285 1 0 $X=120710 $Y=109715
X1196 22 22 22 2 1 ne3i_6_CDNS_7246548160536 $T=128170 100985 0 0 $X=124110 $Y=96535
X1197 22 22 22 2 1 ne3i_6_CDNS_7246548160536 $T=128170 124285 1 0 $X=124110 $Y=109715
X1198 1 1 1 ne3_CDNS_7246548160537 $T=11530 16320 0 0 $X=10730 $Y=15920
X1199 1 1 1 ne3_CDNS_7246548160537 $T=11530 38460 1 0 $X=10730 $Y=27890
X1200 1 13 21 ne3_CDNS_7246548160537 $T=14770 16320 0 0 $X=13970 $Y=15920
X1201 1 13 13 ne3_CDNS_7246548160537 $T=14770 38460 1 0 $X=13970 $Y=27890
X1202 1 13 14 ne3_CDNS_7246548160537 $T=18010 16320 0 0 $X=17210 $Y=15920
X1203 1 13 21 ne3_CDNS_7246548160537 $T=18010 38460 1 0 $X=17210 $Y=27890
X1204 1 13 13 ne3_CDNS_7246548160537 $T=21250 16320 0 0 $X=20450 $Y=15920
X1205 1 13 14 ne3_CDNS_7246548160537 $T=21250 38460 1 0 $X=20450 $Y=27890
X1206 1 13 21 ne3_CDNS_7246548160537 $T=24490 16320 0 0 $X=23690 $Y=15920
X1207 1 13 13 ne3_CDNS_7246548160537 $T=24490 38460 1 0 $X=23690 $Y=27890
X1208 1 13 14 ne3_CDNS_7246548160537 $T=27730 16320 0 0 $X=26930 $Y=15920
X1209 1 13 21 ne3_CDNS_7246548160537 $T=27730 38460 1 0 $X=26930 $Y=27890
X1210 1 13 13 ne3_CDNS_7246548160537 $T=30970 16320 0 0 $X=30170 $Y=15920
X1211 1 13 14 ne3_CDNS_7246548160537 $T=30970 38460 1 0 $X=30170 $Y=27890
X1212 1 13 21 ne3_CDNS_7246548160537 $T=34210 16320 0 0 $X=33410 $Y=15920
X1213 1 13 13 ne3_CDNS_7246548160537 $T=34210 38460 1 0 $X=33410 $Y=27890
X1214 1 13 14 ne3_CDNS_7246548160537 $T=37450 16320 0 0 $X=36650 $Y=15920
X1215 1 13 21 ne3_CDNS_7246548160537 $T=37450 38460 1 0 $X=36650 $Y=27890
X1216 1 13 13 ne3_CDNS_7246548160537 $T=40690 16320 0 0 $X=39890 $Y=15920
X1217 1 13 14 ne3_CDNS_7246548160537 $T=40690 38460 1 0 $X=39890 $Y=27890
X1218 1 13 21 ne3_CDNS_7246548160537 $T=43930 16320 0 0 $X=43130 $Y=15920
X1219 1 13 13 ne3_CDNS_7246548160537 $T=43930 38460 1 0 $X=43130 $Y=27890
X1220 1 13 14 ne3_CDNS_7246548160537 $T=47170 16320 0 0 $X=46370 $Y=15920
X1221 1 13 21 ne3_CDNS_7246548160537 $T=47170 38460 1 0 $X=46370 $Y=27890
X1222 1 13 13 ne3_CDNS_7246548160537 $T=50410 16320 0 0 $X=49610 $Y=15920
X1223 1 13 14 ne3_CDNS_7246548160537 $T=50410 38460 1 0 $X=49610 $Y=27890
X1224 1 1 1 ne3_CDNS_7246548160537 $T=53650 16320 0 0 $X=52850 $Y=15920
X1225 1 1 1 ne3_CDNS_7246548160537 $T=53650 38460 1 0 $X=52850 $Y=27890
X1226 2 1 pe3_CDNS_7246548160538 $T=205435 52315 1 0 $X=203925 $Y=49285
X1227 2 1 pe3_CDNS_7246548160538 $T=205435 175915 1 0 $X=203925 $Y=172885
X1228 2 1 pe3_CDNS_7246548160538 $T=216675 52315 1 0 $X=215165 $Y=49285
X1229 2 1 pe3_CDNS_7246548160538 $T=216675 175915 1 0 $X=215165 $Y=172885
X1230 2 1 pe3_CDNS_7246548160538 $T=227915 52315 1 0 $X=226405 $Y=49285
X1231 2 1 pe3_CDNS_7246548160538 $T=227915 175915 1 0 $X=226405 $Y=172885
X1232 2 1 pe3_CDNS_7246548160538 $T=239155 52315 1 0 $X=237645 $Y=49285
X1233 2 1 pe3_CDNS_7246548160538 $T=239155 175915 1 0 $X=237645 $Y=172885
X1234 2 1 pe3_CDNS_7246548160538 $T=250395 52315 1 0 $X=248885 $Y=49285
X1235 2 1 pe3_CDNS_7246548160538 $T=250395 175915 1 0 $X=248885 $Y=172885
X1236 2 1 pe3_CDNS_7246548160538 $T=261635 52315 1 0 $X=260125 $Y=49285
X1237 2 1 pe3_CDNS_7246548160538 $T=261635 175915 1 0 $X=260125 $Y=172885
X1238 2 1 pe3_CDNS_7246548160538 $T=272875 52315 1 0 $X=271365 $Y=49285
X1239 2 1 pe3_CDNS_7246548160538 $T=272875 175915 1 0 $X=271365 $Y=172885
X1240 2 1 pe3_CDNS_7246548160538 $T=284115 52315 1 0 $X=282605 $Y=49285
X1241 2 1 pe3_CDNS_7246548160538 $T=284115 175915 1 0 $X=282605 $Y=172885
X1242 2 1 pe3_CDNS_7246548160538 $T=295355 52315 1 0 $X=293845 $Y=49285
X1243 2 1 pe3_CDNS_7246548160538 $T=295355 175915 1 0 $X=293845 $Y=172885
X1244 2 1 pe3_CDNS_7246548160538 $T=306595 52315 1 0 $X=305085 $Y=49285
X1245 2 1 pe3_CDNS_7246548160538 $T=306595 175915 1 0 $X=305085 $Y=172885
X1246 2 1 pe3_CDNS_7246548160538 $T=317835 52315 1 0 $X=316325 $Y=49285
X1247 2 1 pe3_CDNS_7246548160538 $T=317835 175915 1 0 $X=316325 $Y=172885
X1248 2 1 pe3_CDNS_7246548160538 $T=329075 52315 1 0 $X=327565 $Y=49285
X1249 2 1 pe3_CDNS_7246548160538 $T=329075 175915 1 0 $X=327565 $Y=172885
X1250 2 1 pe3_CDNS_7246548160538 $T=340315 52315 1 0 $X=338805 $Y=49285
X1251 2 1 pe3_CDNS_7246548160538 $T=340315 175915 1 0 $X=338805 $Y=172885
X1252 2 1 pe3_CDNS_7246548160538 $T=351555 52315 1 0 $X=350045 $Y=49285
X1253 2 1 pe3_CDNS_7246548160538 $T=351555 175915 1 0 $X=350045 $Y=172885
X1254 2 1 pe3_CDNS_7246548160538 $T=362795 52315 1 0 $X=361285 $Y=49285
X1255 2 1 pe3_CDNS_7246548160538 $T=362795 175915 1 0 $X=361285 $Y=172885
X1256 1 25 13 ne3_CDNS_7246548160539 $T=96785 56345 0 0 $X=95985 $Y=55765
X1257 1 25 5 ne3_CDNS_7246548160539 $T=102390 56345 0 0 $X=101590 $Y=55765
X1258 2 2 2 17 16 16 17 1 MASCO__A15 $T=54830 160530 0 0 $X=54830 $Y=160530
X1259 16 16 2 17 16 16 17 1 MASCO__A15 $T=99790 160530 0 0 $X=99790 $Y=160530
X1260 2 2 2 26 17 27 27 1 MASCO__A15 $T=203925 60085 0 0 $X=203925 $Y=60085
X1261 2 2 2 26 17 27 28 1 MASCO__A15 $T=203925 78885 0 0 $X=203925 $Y=78885
X1262 2 2 2 26 17 27 28 1 MASCO__A15 $T=203925 97685 0 0 $X=203925 $Y=97685
X1263 2 2 2 26 17 27 28 1 MASCO__A15 $T=203925 116485 0 0 $X=203925 $Y=116485
X1264 2 2 2 26 17 27 28 1 MASCO__A15 $T=203925 135285 0 0 $X=203925 $Y=135285
X1265 2 2 2 26 17 26 26 1 MASCO__A15 $T=203925 154085 0 0 $X=203925 $Y=154085
X1266 27 17 2 27 17 30 26 1 MASCO__A15 $T=248885 60085 0 0 $X=248885 $Y=60085
X1267 30 17 2 31 17 31 30 1 MASCO__A15 $T=248885 78885 0 0 $X=248885 $Y=78885
X1268 29 17 2 30 17 24 30 1 MASCO__A15 $T=248885 97685 0 0 $X=248885 $Y=97685
X1269 30 17 2 29 17 30 28 1 MASCO__A15 $T=248885 116485 0 0 $X=248885 $Y=116485
X1270 30 17 2 31 17 31 30 1 MASCO__A15 $T=248885 135285 0 0 $X=248885 $Y=135285
X1271 26 17 2 26 17 27 27 1 MASCO__A15 $T=248885 154085 0 0 $X=248885 $Y=154085
X1272 26 17 2 2 2 2 2 1 MASCO__A15 $T=293845 60085 0 0 $X=293845 $Y=60085
X1273 28 17 2 27 17 26 26 1 MASCO__A15 $T=293845 78885 0 0 $X=293845 $Y=78885
X1274 28 17 2 27 17 26 26 1 MASCO__A15 $T=293845 97685 0 0 $X=293845 $Y=97685
X1275 27 17 2 27 17 26 26 1 MASCO__A15 $T=293845 116485 0 0 $X=293845 $Y=116485
X1276 28 17 2 27 17 26 26 1 MASCO__A15 $T=293845 135285 0 0 $X=293845 $Y=135285
X1277 27 17 2 30 17 26 26 1 MASCO__A15 $T=293845 154085 0 0 $X=293845 $Y=154085
D0 1 2 p_dnw AREA=7.95604e-10 PJ=0.00014876 perimeter=0.00014876 $X=8500 $Y=140710 $dt=6
D1 1 2 p_dnw AREA=2.14716e-09 PJ=0.0003306 perimeter=0.0003306 $X=48630 $Y=140710 $dt=6
D2 1 2 p_dnw AREA=3.11448e-11 PJ=3.188e-05 perimeter=3.188e-05 $X=88435 $Y=59745 $dt=6
D3 1 18 p_dnw AREA=1.97548e-10 PJ=8.944e-05 perimeter=8.944e-05 $X=151005 $Y=72505 $dt=6
D4 1 19 p_dnw AREA=1.97548e-10 PJ=8.944e-05 perimeter=8.944e-05 $X=151005 $Y=93985 $dt=6
D5 1 20 p_dnw AREA=1.97548e-10 PJ=8.944e-05 perimeter=8.944e-05 $X=151005 $Y=114935 $dt=6
D6 1 2 p_dnw AREA=1.47356e-08 PJ=0.0006944 perimeter=0.0006944 $X=181765 $Y=46865 $dt=6
D7 1 2 p_dnw AREA=1.65707e-09 PJ=0.00035483 perimeter=0.00035483 $X=220785 $Y=22870 $dt=6
D8 1 2 p_dnw AREA=6.02548e-10 PJ=0.00014223 perimeter=0.00014223 $X=303405 $Y=4665 $dt=6
D9 1 2 p_ddnw AREA=1.72778e-09 PJ=0.0002104 perimeter=0.0002104 $X=65040 $Y=95265 $dt=7
D10 22 2 p_dipdnwmv AREA=9.7703e-10 PJ=0.0001796 perimeter=0.0001796 $X=68890 $Y=99115 $dt=8
D11 1 2 p_dnw3 AREA=2.92576e-10 PJ=0 perimeter=0 $X=14200 $Y=147550 $dt=9
D12 1 2 p_dnw3 AREA=2.92576e-10 PJ=0 perimeter=0 $X=14200 $Y=160530 $dt=9
D13 1 2 p_dnw3 AREA=1.37701e-09 PJ=0 perimeter=0 $X=54830 $Y=147550 $dt=9
D14 1 2 p_dnw3 AREA=1.37701e-09 PJ=0 perimeter=0 $X=54830 $Y=160530 $dt=9
D15 1 2 p_dnw3 AREA=2.67592e-11 PJ=0 perimeter=0 $X=89575 $Y=60885 $dt=9
D16 1 18 p_dnw3 AREA=2.77621e-10 PJ=0 perimeter=0 $X=153165 $Y=75665 $dt=9
D17 1 19 p_dnw3 AREA=2.77621e-10 PJ=0 perimeter=0 $X=153165 $Y=97145 $dt=9
D18 1 20 p_dnw3 AREA=2.77621e-10 PJ=0 perimeter=0 $X=153165 $Y=118095 $dt=9
D19 1 2 p_dnw3 AREA=6.91743e-10 PJ=0 perimeter=0 $X=203925 $Y=49285 $dt=9
D20 1 2 p_dnw3 AREA=2.05478e-09 PJ=0 perimeter=0 $X=203925 $Y=60085 $dt=9
D21 1 2 p_dnw3 AREA=2.05478e-09 PJ=0 perimeter=0 $X=203925 $Y=78885 $dt=9
D22 1 2 p_dnw3 AREA=2.05478e-09 PJ=0 perimeter=0 $X=203925 $Y=97685 $dt=9
D23 1 2 p_dnw3 AREA=2.05478e-09 PJ=0 perimeter=0 $X=203925 $Y=116485 $dt=9
D24 1 2 p_dnw3 AREA=2.05478e-09 PJ=0 perimeter=0 $X=203925 $Y=135285 $dt=9
D25 1 2 p_dnw3 AREA=2.05478e-09 PJ=0 perimeter=0 $X=203925 $Y=154085 $dt=9
D26 1 2 p_dnw3 AREA=6.91743e-10 PJ=0 perimeter=0 $X=203925 $Y=172885 $dt=9
D27 1 2 p_dnw3 AREA=2.15633e-10 PJ=0 perimeter=0 $X=222425 $Y=25290 $dt=9
D28 1 2 p_dnw3 AREA=6.24226e-10 PJ=0 perimeter=0 $X=245245 $Y=25290 $dt=9
D29 1 2 p_dnw3 AREA=3.27067e-10 PJ=0 perimeter=0 $X=301060 $Y=25290 $dt=9
D30 1 2 p_dnw3 AREA=5.13756e-11 PJ=0 perimeter=0 $X=305565 $Y=6305 $dt=9
D31 1 2 p_dnw3 AREA=5.13756e-11 PJ=0 perimeter=0 $X=314825 $Y=6305 $dt=9
D32 1 2 p_dnw3 AREA=5.13756e-11 PJ=0 perimeter=0 $X=324085 $Y=6305 $dt=9
D33 1 2 p_dnw3 AREA=1.78488e-10 PJ=0 perimeter=0 $X=331825 $Y=25290 $dt=9
D34 1 2 p_dnw3 AREA=5.13756e-11 PJ=0 perimeter=0 $X=333345 $Y=6305 $dt=9
D35 1 2 p_dnw3 AREA=5.13756e-11 PJ=0 perimeter=0 $X=342605 $Y=6305 $dt=9
D36 1 2 p_dnw3 AREA=1.04198e-10 PJ=0 perimeter=0 $X=350290 $Y=25290 $dt=9
D37 1 2 p_dnw3 AREA=5.13756e-11 PJ=0 perimeter=0 $X=351865 $Y=6305 $dt=9
D38 1 2 p_dnw3 AREA=6.70536e-11 PJ=0 perimeter=0 $X=362625 $Y=25290 $dt=9
D39 1 2 p_dnw3 AREA=4.84812e-11 PJ=0 perimeter=0 $X=372000 $Y=25290 $dt=9
.ends dac6b_amp_n2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pulse_generator                                 *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pulse_generator 13 7 12 19 18 17 16 15 14 3
+ 8 5 10 4 6 11 2 9
** N=19 EP=18 FDC=594
X0 1 VIA3_C_CDNS_724654816050 $T=510235 23750 0 0 $X=509485 $Y=23000
X1 2 VIA3_C_CDNS_724654816051 $T=75160 135625 0 0 $X=74410 $Y=135395
X2 3 VIA3_C_CDNS_724654816051 $T=79660 101100 0 0 $X=78910 $Y=100870
X3 2 VIA3_C_CDNS_724654816052 $T=74075 135625 0 0 $X=73935 $Y=135375
X4 3 VIA3_C_CDNS_724654816052 $T=78295 101100 0 0 $X=78155 $Y=100850
X5 3 VIA3_C_CDNS_724654816053 $T=424330 102600 0 0 $X=423580 $Y=102110
X6 4 VIA3_C_CDNS_724654816053 $T=428475 102625 0 0 $X=427725 $Y=102135
X7 5 6 3 7 4 1 8 9 10 11
+ 12 current_source_gm_10_en_r $T=412080 18790 0 0 $X=416015 $Y=22610
X8 5 6 mosvc3_CDNS_7246548160521 $T=21090 101820 0 0 $X=20290 $Y=101390
X9 5 6 mosvc3_CDNS_7246548160521 $T=21090 154080 1 0 $X=20290 $Y=128460
X10 5 6 mosvc3_CDNS_7246548160521 $T=44090 101820 0 0 $X=43290 $Y=101390
X11 5 6 mosvc3_CDNS_7246548160521 $T=44090 154080 1 0 $X=43290 $Y=128460
X12 5 6 mosvc3_CDNS_7246548160522 $T=422175 183935 0 0 $X=421375 $Y=183505
X13 5 6 mosvc3_CDNS_7246548160522 $T=445175 183935 0 0 $X=444375 $Y=183505
X14 5 6 mosvc3_CDNS_7246548160522 $T=468175 183935 0 0 $X=467375 $Y=183505
X15 5 6 mosvc3_CDNS_7246548160522 $T=491175 183935 0 0 $X=490375 $Y=183505
X16 5 6 mosvc3_CDNS_7246548160522 $T=514175 183935 0 0 $X=513375 $Y=183505
X17 5 6 mosvc3_CDNS_7246548160522 $T=537175 183935 0 0 $X=536375 $Y=183505
X18 5 6 mosvc3_CDNS_7246548160522 $T=560175 183935 0 0 $X=559375 $Y=183505
X19 5 6 mosvc3_CDNS_7246548160522 $T=583175 183935 0 0 $X=582375 $Y=183505
X20 5 6 13 3 1 2 14 15 16 17
+ 18 19 dac6b_amp_n2 $T=14140 23390 0 0 $X=16780 $Y=24625
R0 5 9 5 $[s_res] $X=675360 $Y=22605 $dt=5
.ends pulse_generator
