* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : constant_gm                                  *
* Netlisted  : Mon Aug 26 08:12:02 2024                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(ne3) nem ndiff(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 1 MP(pe3) pem pdiff(D) p1trm(G) pdiff(S) nwtrm(B)
*.DEVTMPLT 2 NE3I_6() nemi_6 ndiff(D) p1trm(G) ndiff(S) pwitrm(B) dnwtrm(NW) bulk(SB)
*.DEVTMPLT 3 D(p_dnw) p_dnw bulk(POS) nwtrm(NEG)
*.DEVTMPLT 4 D(p_ddnw) p_ddnw bulk(POS) dnwtrm(NEG)
*.DEVTMPLT 5 D(p_dipdnwmv) p_dipwmv pwitrm(POS) dnwtrm(NEG)
*.DEVTMPLT 6 D(p_dnw3) p_dnwm bulk(POS) nwtrm(NEG)
*.DEVTMPLT 7 R(rpp1k1_3) rpp1k1_n p1trm(POS) p1trm(NEG) nwtrm(SUB)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724652717070                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724652717070 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724652717070

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724652717072                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724652717072 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724652717072

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724652717073                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724652717073 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724652717073

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_724652717077                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_724652717077 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_724652717077

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_724652717078                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_724652717078 1
*.DEVICECLIMB
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_724652717078

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724652717079                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724652717079 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724652717079

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246527170711                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246527170711 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246527170711

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246527170712                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246527170712 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246527170712

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246527170713                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246527170713 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246527170713

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246527170718                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246527170718 1 2
*.DEVICECLIMB
** N=2 EP=2 FDC=0
.ends VIA2_C_CDNS_7246527170718

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246527170719                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246527170719 1 2
** N=2 EP=2 FDC=0
.ends VIA2_C_CDNS_7246527170719

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3i_6_CDNS_724652717070                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3i_6_CDNS_724652717070 1 2 3
** N=3 EP=3 FDC=4
X0 1 3 3 1 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=4.8e-12 ps=1.054e-05 pd=2.096e-05 $X=0 $Y=0 $dt=2
X1 3 3 1 1 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=4.8e-12 ad=2.7e-12 ps=2.096e-05 pd=1.054e-05 $X=3040 $Y=0 $dt=2
D2 1 2 p_ddnw AREA=3.07331e-10 PJ=7.576e-05 perimeter=7.576e-05 $X=-6110 $Y=-4940 $dt=4
D3 1 2 p_dipdnwmv AREA=7.49452e-11 PJ=4.496e-05 perimeter=4.496e-05 $X=-2260 $Y=-1090 $dt=5
.ends ne3i_6_CDNS_724652717070

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724652717071                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724652717071 1 2 3
** N=3 EP=3 FDC=2
M0 2 2 1 1 pe3 L=1e-05 W=2e-06 AD=9.6e-13 AS=9.6e-13 PD=4.96e-06 PS=4.96e-06 $X=0 $Y=0 $dt=1
D1 3 1 p_dnw3 AREA=4.57434e-11 PJ=3.138e-05 perimeter=3.138e-05 $X=-910 $Y=-1440 $dt=6
.ends pe3_CDNS_724652717071

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724652717072                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724652717072 1 2 3 4
** N=4 EP=4 FDC=2
M0 3 2 1 4 ne3 L=2.5e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
M1 1 2 3 4 ne3 L=2.5e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=3040 $Y=0 $dt=0
.ends ne3_CDNS_724652717072

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724652717073                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724652717073 1 2 3 4 5
** N=5 EP=5 FDC=3
M0 3 2 1 4 pe3 L=2.5e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=2.5e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=3040 $Y=0 $dt=1
D2 5 4 p_dnw3 AREA=1.03234e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=6
.ends pe3_CDNS_724652717073

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724652717074                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724652717074 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 3 2 1 4 pe3 L=2.5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
D1 5 4 p_dnw3 AREA=6.65712e-11 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=6
.ends pe3_CDNS_724652717074

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724652717075                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724652717075 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
M0 3 2 1 1 pe3 L=2.5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_724652717075

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3i_6_CDNS_724652717076                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3i_6_CDNS_724652717076 1 2 3 4 5
** N=5 EP=5 FDC=10
X0 3 4 5 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=4.8e-12 ps=1.054e-05 pd=2.096e-05 $X=0 $Y=0 $dt=2
X1 5 4 3 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=2.7e-12 ps=1.054e-05 pd=1.054e-05 $X=3040 $Y=0 $dt=2
X2 3 4 5 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=2.7e-12 ps=1.054e-05 pd=1.054e-05 $X=6080 $Y=0 $dt=2
X3 5 4 3 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=2.7e-12 ps=1.054e-05 pd=1.054e-05 $X=9120 $Y=0 $dt=2
X4 3 4 5 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=2.7e-12 ps=1.054e-05 pd=1.054e-05 $X=12160 $Y=0 $dt=2
X5 5 4 3 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=2.7e-12 ps=1.054e-05 pd=1.054e-05 $X=15200 $Y=0 $dt=2
X6 3 4 5 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=2.7e-12 ps=1.054e-05 pd=1.054e-05 $X=18240 $Y=0 $dt=2
X7 5 4 3 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=4.8e-12 ad=2.7e-12 ps=2.096e-05 pd=1.054e-05 $X=21280 $Y=0 $dt=2
D8 1 2 p_ddnw AREA=5.2432e-10 PJ=0.00011224 perimeter=0.00011224 $X=-6110 $Y=-4940 $dt=4
D9 3 2 p_dipdnwmv AREA=1.51486e-10 PJ=8.144e-05 perimeter=8.144e-05 $X=-2260 $Y=-1090 $dt=5
.ends ne3i_6_CDNS_724652717076

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_724652717077                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_724652717077 1 2 3
*.DEVICECLIMB
** N=3 EP=3 FDC=1
R0 2 1 L=0.0002878 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=7
.ends rpp1k1_3_CDNS_724652717077

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: constant_gm                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt constant_gm 13 9 11 16 14
** N=16 EP=5 FDC=56
X0 1 VIA1_C_CDNS_724652717070 $T=11390 57075 0 0 $X=10990 $Y=56625
X1 2 VIA1_C_CDNS_724652717070 $T=14430 55795 0 0 $X=14030 $Y=55345
X2 1 VIA1_C_CDNS_724652717070 $T=17470 57075 0 0 $X=17070 $Y=56625
X3 3 VIA1_C_CDNS_724652717070 $T=21540 55655 0 0 $X=21140 $Y=55205
X4 4 VIA1_C_CDNS_724652717070 $T=24580 56935 0 0 $X=24180 $Y=56485
X5 5 VIA1_C_CDNS_724652717070 $T=25190 37045 0 0 $X=24790 $Y=36595
X6 6 VIA1_C_CDNS_724652717070 $T=25275 95030 0 0 $X=24875 $Y=94580
X7 6 VIA1_C_CDNS_724652717070 $T=25275 114390 0 0 $X=24875 $Y=113940
X8 3 VIA1_C_CDNS_724652717070 $T=27620 55655 0 0 $X=27220 $Y=55205
X9 2 VIA1_C_CDNS_724652717070 $T=28230 38325 0 0 $X=27830 $Y=37875
X10 1 VIA1_C_CDNS_724652717070 $T=29015 111830 0 0 $X=28615 $Y=111380
X11 5 VIA1_C_CDNS_724652717070 $T=31270 37045 0 0 $X=30870 $Y=36595
X12 7 VIA1_C_CDNS_724652717070 $T=32295 55655 0 0 $X=31895 $Y=55205
X13 1 VIA1_C_CDNS_724652717070 $T=32755 92470 0 0 $X=32355 $Y=92020
X14 8 VIA1_C_CDNS_724652717070 $T=34520 37045 0 0 $X=34120 $Y=36595
X15 9 VIA1_C_CDNS_724652717070 $T=35335 56935 0 0 $X=34935 $Y=56485
X16 7 VIA1_C_CDNS_724652717070 $T=36495 93750 0 0 $X=36095 $Y=93300
X17 7 VIA1_C_CDNS_724652717070 $T=36495 113110 0 0 $X=36095 $Y=112660
X18 4 VIA1_C_CDNS_724652717070 $T=37560 38325 0 0 $X=37160 $Y=37875
X19 7 VIA1_C_CDNS_724652717070 $T=38375 55655 0 0 $X=37975 $Y=55205
X20 10 VIA1_C_CDNS_724652717070 $T=40235 115670 0 0 $X=39835 $Y=115220
X21 8 VIA1_C_CDNS_724652717070 $T=40600 37045 0 0 $X=40200 $Y=36595
X22 6 VIA1_C_CDNS_724652717070 $T=43110 55655 0 0 $X=42710 $Y=55205
X23 11 VIA1_C_CDNS_724652717070 $T=46150 56935 0 0 $X=45750 $Y=56485
X24 6 VIA1_C_CDNS_724652717070 $T=49190 55655 0 0 $X=48790 $Y=55205
X25 3 VIA1_C_CDNS_724652717072 $T=23755 75790 0 0 $X=23615 $Y=75340
X26 3 VIA1_C_CDNS_724652717072 $T=23755 91190 0 0 $X=23615 $Y=90740
X27 3 VIA1_C_CDNS_724652717072 $T=27495 75790 0 0 $X=27355 $Y=75340
X28 3 VIA1_C_CDNS_724652717072 $T=27495 91190 0 0 $X=27355 $Y=90740
X29 3 VIA1_C_CDNS_724652717072 $T=31235 75790 0 0 $X=31095 $Y=75340
X30 3 VIA1_C_CDNS_724652717072 $T=31235 91190 0 0 $X=31095 $Y=90740
X31 3 VIA1_C_CDNS_724652717072 $T=34975 75790 0 0 $X=34835 $Y=75340
X32 3 VIA1_C_CDNS_724652717072 $T=34975 91190 0 0 $X=34835 $Y=90740
X33 3 VIA1_C_CDNS_724652717072 $T=38715 91190 0 0 $X=38575 $Y=90740
X34 12 VIA1_C_CDNS_724652717073 $T=64765 41965 0 0 $X=62975 $Y=41475
X35 13 VIA1_C_CDNS_724652717073 $T=77600 41965 0 0 $X=75810 $Y=41475
X36 13 VIA1_C_CDNS_724652717073 $T=77650 33280 0 0 $X=75860 $Y=32790
X37 9 VIA2_C_CDNS_724652717077 $T=35335 56935 0 0 $X=33805 $Y=56445
X38 8 VIA2_C_CDNS_724652717077 $T=36610 37055 0 0 $X=35080 $Y=36565
X39 11 VIA2_C_CDNS_724652717077 $T=46150 56935 0 0 $X=44620 $Y=56445
X40 14 VIA2_C_CDNS_724652717078 $T=16225 89660 0 0 $X=15515 $Y=89000
X41 14 VIA2_C_CDNS_724652717078 $T=16225 109020 0 0 $X=15515 $Y=108360
X42 14 VIA2_C_CDNS_724652717078 $T=46245 89660 0 0 $X=45535 $Y=89000
X43 14 VIA2_C_CDNS_724652717078 $T=46245 109020 0 0 $X=45535 $Y=108360
X44 14 VIA1_C_CDNS_724652717079 $T=18495 89660 0 0 $X=18355 $Y=88950
X45 14 VIA1_C_CDNS_724652717079 $T=18495 109020 0 0 $X=18355 $Y=108310
X46 14 VIA1_C_CDNS_724652717079 $T=21535 89660 0 0 $X=21395 $Y=88950
X47 14 VIA1_C_CDNS_724652717079 $T=21535 109020 0 0 $X=21395 $Y=108310
X48 14 VIA1_C_CDNS_724652717079 $T=22235 89660 0 0 $X=22095 $Y=88950
X49 14 VIA1_C_CDNS_724652717079 $T=22235 109020 0 0 $X=22095 $Y=108310
X50 14 VIA1_C_CDNS_724652717079 $T=25975 89660 0 0 $X=25835 $Y=88950
X51 14 VIA1_C_CDNS_724652717079 $T=25975 109020 0 0 $X=25835 $Y=108310
X52 14 VIA1_C_CDNS_724652717079 $T=29715 89660 0 0 $X=29575 $Y=88950
X53 14 VIA1_C_CDNS_724652717079 $T=29715 109020 0 0 $X=29575 $Y=108310
X54 14 VIA1_C_CDNS_724652717079 $T=33455 89660 0 0 $X=33315 $Y=88950
X55 14 VIA1_C_CDNS_724652717079 $T=33455 109020 0 0 $X=33315 $Y=108310
X56 14 VIA1_C_CDNS_724652717079 $T=37195 89660 0 0 $X=37055 $Y=88950
X57 14 VIA1_C_CDNS_724652717079 $T=37195 109020 0 0 $X=37055 $Y=108310
X58 14 VIA1_C_CDNS_724652717079 $T=40235 89660 0 0 $X=40095 $Y=88950
X59 14 VIA1_C_CDNS_724652717079 $T=40935 89660 0 0 $X=40795 $Y=88950
X60 14 VIA1_C_CDNS_724652717079 $T=40935 109020 0 0 $X=40795 $Y=108310
X61 14 VIA1_C_CDNS_724652717079 $T=43975 89660 0 0 $X=43835 $Y=88950
X62 14 VIA1_C_CDNS_724652717079 $T=43975 109020 0 0 $X=43835 $Y=108310
X63 1 VIA2_C_CDNS_7246527170711 $T=14445 92470 0 0 $X=13735 $Y=92070
X64 1 VIA2_C_CDNS_7246527170711 $T=14445 111830 0 0 $X=13735 $Y=111430
X65 3 VIA2_C_CDNS_7246527170711 $T=48025 75790 0 0 $X=47315 $Y=75390
X66 3 VIA2_C_CDNS_7246527170711 $T=48025 91190 0 0 $X=47315 $Y=90790
X67 3 VIA2_C_CDNS_7246527170711 $T=48025 110550 0 0 $X=47315 $Y=110150
X68 7 VIA2_C_CDNS_7246527170711 $T=49805 93750 0 0 $X=49095 $Y=93350
X69 7 VIA2_C_CDNS_7246527170711 $T=49805 113110 0 0 $X=49095 $Y=112710
X70 6 VIA2_C_CDNS_7246527170711 $T=51585 95030 0 0 $X=50875 $Y=94630
X71 6 VIA2_C_CDNS_7246527170711 $T=51585 114390 0 0 $X=50875 $Y=113990
X72 10 VIA2_C_CDNS_7246527170711 $T=53365 115670 0 0 $X=52655 $Y=115270
X73 3 VIA1_C_CDNS_7246527170712 $T=29015 91190 0 0 $X=28045 $Y=91050
X74 3 VIA1_C_CDNS_7246527170712 $T=32755 110550 0 0 $X=31785 $Y=110410
X75 4 VIA1_C_CDNS_7246527170713 $T=12910 70305 0 0 $X=11990 $Y=70115
X76 4 VIA1_C_CDNS_7246527170713 $T=15950 70305 0 0 $X=15030 $Y=70115
X77 4 VIA1_C_CDNS_7246527170713 $T=23060 70305 0 0 $X=22140 $Y=70115
X78 4 VIA1_C_CDNS_7246527170713 $T=26100 70305 0 0 $X=25180 $Y=70115
X79 2 VIA1_C_CDNS_7246527170713 $T=26710 50605 0 0 $X=25790 $Y=50415
X80 2 VIA1_C_CDNS_7246527170713 $T=29750 50605 0 0 $X=28830 $Y=50415
X81 4 VIA1_C_CDNS_7246527170713 $T=33815 70305 0 0 $X=32895 $Y=70115
X82 2 VIA1_C_CDNS_7246527170713 $T=36040 50605 0 0 $X=35120 $Y=50415
X83 4 VIA1_C_CDNS_7246527170713 $T=36855 70305 0 0 $X=35935 $Y=70115
X84 2 VIA1_C_CDNS_7246527170713 $T=39080 50605 0 0 $X=38160 $Y=50415
X85 4 VIA1_C_CDNS_7246527170713 $T=44630 70305 0 0 $X=43710 $Y=70115
X86 4 VIA1_C_CDNS_7246527170713 $T=47670 70305 0 0 $X=46750 $Y=70115
X87 1 14 VIA2_C_CDNS_7246527170718 $T=19200 68420 0 0 $X=18450 $Y=67760
X88 3 14 VIA2_C_CDNS_7246527170718 $T=29865 68705 0 0 $X=29115 $Y=68045
X89 7 14 VIA2_C_CDNS_7246527170718 $T=40615 68490 0 0 $X=39865 $Y=67830
X90 14 13 VIA2_C_CDNS_7246527170719 $T=16225 120015 0 0 $X=14695 $Y=118485
X91 14 13 VIA2_C_CDNS_7246527170719 $T=46240 119870 0 0 $X=44710 $Y=118340
X92 13 14 5 ne3i_6_CDNS_724652717070 $T=18020 14875 0 0 $X=7250 $Y=5275
X93 15 2 13 pe3_CDNS_724652717071 $T=10155 41775 0 0 $X=8645 $Y=39735
X94 4 15 13 pe3_CDNS_724652717071 $T=20155 47905 1 180 $X=8645 $Y=45865
X95 5 2 2 13 ne3_CDNS_724652717072 $T=25460 39505 0 0 $X=24660 $Y=39105
X96 8 2 4 13 ne3_CDNS_724652717072 $T=34790 39505 0 0 $X=33990 $Y=39105
X97 1 4 2 14 13 pe3_CDNS_724652717073 $T=11660 58745 0 0 $X=10150 $Y=57715
X98 3 4 4 14 13 pe3_CDNS_724652717073 $T=21810 58745 0 0 $X=20300 $Y=57715
X99 7 4 9 14 13 pe3_CDNS_724652717073 $T=32565 58745 0 0 $X=31055 $Y=57715
X100 6 4 11 14 13 pe3_CDNS_724652717073 $T=43380 58745 0 0 $X=41870 $Y=57715
X101 10 4 16 14 13 pe3_CDNS_724652717074 $T=53845 58745 0 0 $X=52335 $Y=57715
X102 14 14 14 13 pe3_CDNS_724652717075 $T=18765 87600 1 0 $X=17255 $Y=76570
X103 14 14 14 13 pe3_CDNS_724652717075 $T=18765 106960 1 0 $X=17255 $Y=95930
X104 14 3 6 13 pe3_CDNS_724652717075 $T=22505 87600 1 0 $X=20995 $Y=76570
X105 14 3 6 13 pe3_CDNS_724652717075 $T=22505 106960 1 0 $X=20995 $Y=95930
X106 14 3 3 13 pe3_CDNS_724652717075 $T=26245 87600 1 0 $X=24735 $Y=76570
X107 14 3 1 13 pe3_CDNS_724652717075 $T=26245 106960 1 0 $X=24735 $Y=95930
X108 14 3 1 13 pe3_CDNS_724652717075 $T=29985 87600 1 0 $X=28475 $Y=76570
X109 14 3 3 13 pe3_CDNS_724652717075 $T=29985 106960 1 0 $X=28475 $Y=95930
X110 14 3 7 13 pe3_CDNS_724652717075 $T=33725 87600 1 0 $X=32215 $Y=76570
X111 14 3 7 13 pe3_CDNS_724652717075 $T=33725 106960 1 0 $X=32215 $Y=95930
X112 14 14 14 13 pe3_CDNS_724652717075 $T=37465 87600 1 0 $X=35955 $Y=76570
X113 14 3 10 13 pe3_CDNS_724652717075 $T=37465 106960 1 0 $X=35955 $Y=95930
X114 14 14 14 13 pe3_CDNS_724652717075 $T=41205 87600 1 0 $X=39695 $Y=76570
X115 14 14 14 13 pe3_CDNS_724652717075 $T=41205 106960 1 0 $X=39695 $Y=95930
X116 13 14 12 5 8 ne3i_6_CDNS_724652717076 $T=48275 14875 0 0 $X=37505 $Y=5275
X117 13 12 14 rpp1k1_3_CDNS_724652717077 $T=62765 46455 1 90 $X=62545 $Y=41295
D0 13 14 p_dnw AREA=4.77568e-10 PJ=0.00014131 perimeter=0.00014131 $X=7700 $Y=53605 $dt=3
D1 13 14 p_dnw AREA=1.16854e-09 PJ=0.00017172 perimeter=0.00017172 $X=12555 $Y=74150 $dt=3
D2 13 14 p_dnw AREA=1.48411e-09 PJ=0.00019385 perimeter=0.00019385 $X=61625 $Y=40375 $dt=3
D3 13 14 p_dnw3 AREA=3.37198e-10 PJ=0 perimeter=0 $X=17255 $Y=76570 $dt=6
D4 13 14 p_dnw3 AREA=3.37198e-10 PJ=0 perimeter=0 $X=17255 $Y=95930 $dt=6
.ends constant_gm
