* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : dac6b_amp_n2                                 *
* Netlisted  : Wed Jun 26 14:49:12 2024                     *
* PVS Version: 23.10-p043 Mon Oct 2 18:09:08 PDT 2023      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(ne3) nem ndiff(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 1 MP(pe3) pem pdiff(D) p1trm(G) pdiff(S) nwtrm(B)
*.DEVTMPLT 2 NE3I_6() nemi_6 ndiff(D) p1trm(G) ndiff(S) pwitrm(B) dnwtrm(NW) bulk(SB)
*.DEVTMPLT 3 D(p_dnw) p_dnw bulk(POS) nwtrm(NEG)
*.DEVTMPLT 4 D(p_ddnw) p_ddnw bulk(POS) dnwtrm(NEG)
*.DEVTMPLT 5 D(p_dipdnwmv) p_dipwmv pwitrm(POS) dnwtrm(NEG)
*.DEVTMPLT 6 D(p_dnw3) p_dnwm bulk(POS) nwtrm(NEG)
*.DEVTMPLT 7 R(rpp1k1_3) rpp1k1_s p1trm(POS) p1trm(NEG) bulk(SUB)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NE3I_6                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NE3I_6 D G S B NW SB
.ends NE3I_6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_719427747080                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_719427747080 1 2 3
*.DEVICECLIMB
** N=4 EP=3 FDC=1
M0 3 2 1 1 pe3 L=1e-05 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_719427747080

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_719427747081                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_719427747081 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
D1 5 4 p_dnw3 AREA=4.84812e-11 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=6
.ends pe3_CDNS_719427747081

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_719427747082                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_719427747082 1 2 3 4 5
** N=5 EP=5 FDC=3
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=1
D2 5 4 p_dnw3 AREA=6.70536e-11 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=6
.ends pe3_CDNS_719427747082

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_719427747083                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_719427747083 1 2 3 4 5
** N=5 EP=5 FDC=5
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=1
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=1
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=1
D4 5 4 p_dnw3 AREA=1.04198e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=6
.ends pe3_CDNS_719427747083

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_719427747084                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_719427747084 1 2 3 4 5
** N=5 EP=5 FDC=9
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=1
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=1
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=1
M4 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=6160 $Y=0 $dt=1
M5 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7700 $Y=0 $dt=1
M6 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=9240 $Y=0 $dt=1
M7 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=10780 $Y=0 $dt=1
D8 5 4 p_dnw3 AREA=1.78488e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=6
.ends pe3_CDNS_719427747084

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_719427747085                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_719427747085 1 2 3 4 5
** N=5 EP=5 FDC=17
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=1
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=1
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=1
M4 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=6160 $Y=0 $dt=1
M5 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7700 $Y=0 $dt=1
M6 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=9240 $Y=0 $dt=1
M7 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10780 $Y=0 $dt=1
M8 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12320 $Y=0 $dt=1
M9 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=13860 $Y=0 $dt=1
M10 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=15400 $Y=0 $dt=1
M11 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=16940 $Y=0 $dt=1
M12 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=18480 $Y=0 $dt=1
M13 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=20020 $Y=0 $dt=1
M14 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=21560 $Y=0 $dt=1
M15 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=23100 $Y=0 $dt=1
D16 5 4 p_dnw3 AREA=3.27067e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=6
.ends pe3_CDNS_719427747085

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_719427747086                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_719427747086 1 2 3 4 5
** N=5 EP=5 FDC=33
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=1
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=1
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=1
M4 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=6160 $Y=0 $dt=1
M5 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7700 $Y=0 $dt=1
M6 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=9240 $Y=0 $dt=1
M7 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10780 $Y=0 $dt=1
M8 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12320 $Y=0 $dt=1
M9 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=13860 $Y=0 $dt=1
M10 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=15400 $Y=0 $dt=1
M11 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=16940 $Y=0 $dt=1
M12 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=18480 $Y=0 $dt=1
M13 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=20020 $Y=0 $dt=1
M14 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=21560 $Y=0 $dt=1
M15 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=23100 $Y=0 $dt=1
M16 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=24640 $Y=0 $dt=1
M17 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=26180 $Y=0 $dt=1
M18 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=27720 $Y=0 $dt=1
M19 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=29260 $Y=0 $dt=1
M20 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=30800 $Y=0 $dt=1
M21 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=32340 $Y=0 $dt=1
M22 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=33880 $Y=0 $dt=1
M23 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=35420 $Y=0 $dt=1
M24 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=36960 $Y=0 $dt=1
M25 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=38500 $Y=0 $dt=1
M26 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=40040 $Y=0 $dt=1
M27 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=41580 $Y=0 $dt=1
M28 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=43120 $Y=0 $dt=1
M29 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=44660 $Y=0 $dt=1
M30 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=46200 $Y=0 $dt=1
M31 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=47740 $Y=0 $dt=1
D32 5 4 p_dnw3 AREA=6.24226e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=6
.ends pe3_CDNS_719427747086

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_719427747087                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_719427747087 1 2
** N=2 EP=2 FDC=1
R0 2 1 L=0.00021702 W=4e-06 $[rpp1k1_3] $SUB=2 $X=-4220 $Y=0 $dt=7
.ends rpp1k1_3_CDNS_719427747087

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_719427747088                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_719427747088 1 2 3 4 5
** N=5 EP=5 FDC=11
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=1
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=1
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=1
M4 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=6160 $Y=0 $dt=1
M5 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7700 $Y=0 $dt=1
M6 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=9240 $Y=0 $dt=1
M7 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10780 $Y=0 $dt=1
M8 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12320 $Y=0 $dt=1
M9 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=13860 $Y=0 $dt=1
D10 5 4 p_dnw3 AREA=2.15633e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=6
.ends pe3_CDNS_719427747088

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_719427747089                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_719427747089 1 2
** N=2 EP=2 FDC=1
R0 2 1 L=0.0008227 W=4e-06 $[rpp1k1_3] $SUB=2 $X=-4220 $Y=0 $dt=7
.ends rpp1k1_3_CDNS_719427747089

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7194277470810                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7194277470810 1 2 3
** N=3 EP=3 FDC=2
M0 2 2 1 1 pe3 L=2e-05 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
D1 3 1 p_dnw3 AREA=2.77621e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=6
.ends pe3_CDNS_7194277470810

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7194277470811                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7194277470811 1 2 3
*.DEVICECLIMB
** N=4 EP=3 FDC=1
M0 3 2 1 1 pe3 L=3e-07 W=6e-06 AD=2.88e-12 AS=2.88e-12 PD=1.296e-05 PS=1.296e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_7194277470811

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7194277470812                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7194277470812 1 2 3 4
** N=4 EP=4 FDC=3
M0 3 2 1 4 pe3 L=3.5e-07 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=3.5e-07 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=890 $Y=0 $dt=1
D2 3 4 p_dnw3 AREA=5.13756e-11 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=6
.ends pe3_CDNS_7194277470812

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7194277470813                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7194277470813 1 2 3 4
** N=4 EP=4 FDC=8
M0 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
M1 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=2540 $Y=0 $dt=0
M2 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=5080 $Y=0 $dt=0
M3 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7620 $Y=0 $dt=0
M4 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10160 $Y=0 $dt=0
M5 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12700 $Y=0 $dt=0
M6 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=15240 $Y=0 $dt=0
M7 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=17780 $Y=0 $dt=0
.ends ne3_CDNS_7194277470813

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7194277470815                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7194277470815 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=2e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
.ends ne3_CDNS_7194277470815

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7194277470816                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7194277470816 1
*.DEVICECLIMB
** N=2 EP=1 FDC=1
M0 1 1 1 1 pe3 L=1e-05 W=2e-06 AD=9.6e-13 AS=9.6e-13 PD=4.96e-06 PS=4.96e-06 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_7194277470816

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7194277470817                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7194277470817 1 2 3
** N=3 EP=3 FDC=4
M0 3 2 1 1 ne3 L=3.5e-07 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
M1 1 2 3 1 ne3 L=3.5e-07 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=890 $Y=0 $dt=0
M2 3 2 1 1 ne3 L=3.5e-07 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1780 $Y=0 $dt=0
M3 1 2 3 1 ne3 L=3.5e-07 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=2670 $Y=0 $dt=0
.ends ne3_CDNS_7194277470817

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7194277470818                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7194277470818 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=3.5e-07 W=2e-06 AD=9.6e-13 AS=9.6e-13 PD=4.96e-06 PS=4.96e-06 $X=0 $Y=0 $dt=0
.ends ne3_CDNS_7194277470818

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A1 1
*.DEVICECLIMB
** N=2 EP=1 FDC=2
X0 1 pe3_CDNS_7194277470816 $T=1510 3030 1 0 $X=0 $Y=0
X1 1 pe3_CDNS_7194277470816 $T=12750 3030 1 0 $X=11240 $Y=0
.ends MASCO__A1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A2 1 2 3 4 5
*.DEVICECLIMB
** N=6 EP=5 FDC=2
X0 1 4 2 pe3_CDNS_719427747080 $T=1510 11030 1 0 $X=0 $Y=0
X1 1 5 3 pe3_CDNS_719427747080 $T=12750 11030 1 0 $X=11240 $Y=0
.ends MASCO__A2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3i_6_CDNS_7194277470814                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3i_6_CDNS_7194277470814 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=1
X0 1 2 3 1 4 5 NE3I_6 w=1e-05 l=2e-06 as=4.8e-12 ad=4.8e-12 ps=2.096e-05 pd=2.096e-05 $X=0 $Y=0 $dt=2
.ends ne3i_6_CDNS_7194277470814

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A3                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A3 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=2
X0 1 3 2 6 7 ne3i_6_CDNS_7194277470814 $T=4060 14570 1 0 $X=0 $Y=0
X1 1 5 4 6 7 ne3i_6_CDNS_7194277470814 $T=7460 14570 1 0 $X=3400 $Y=0
.ends MASCO__A3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A4                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A4 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=2
X0 1 5 4 6 7 ne3i_6_CDNS_7194277470814 $T=4060 4450 0 0 $X=0 $Y=0
X1 1 3 2 6 7 ne3i_6_CDNS_7194277470814 $T=7460 4450 0 0 $X=3400 $Y=0
.ends MASCO__A4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__B5                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__B5 1 2 3 4 5 6 7 8 9 10
+ 11
*.DEVICECLIMB
** N=11 EP=11 FDC=4
X0 1 3 10 5 9 2 11 MASCO__A3 $T=0 13180 0 0 $X=0 $Y=13180
X1 1 6 7 4 8 2 11 MASCO__A4 $T=0 0 0 0 $X=0 $Y=0
.ends MASCO__B5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A6                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A6 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=8 EP=7 FDC=4
X0 1 2 4 7 3 MASCO__A2 $T=0 0 0 0 $X=0 $Y=0
X1 1 5 6 3 3 MASCO__A2 $T=22480 0 0 0 $X=22480 $Y=0
.ends MASCO__A6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: dac6b_amp_n2                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt dac6b_amp_n2 BIAS D0 D1 D2 D3 D4 D5 ENABLE GNDA VDDA
+ VOUT VREF
** N=31 EP=12 FDC=372
X1102 VDDA 4 4 pe3_CDNS_719427747080 $T=15710 148580 0 0 $X=14200 $Y=147550
X1103 VDDA 4 10 pe3_CDNS_719427747080 $T=26950 148580 0 0 $X=25440 $Y=147550
X1104 VDDA VDDA VDDA pe3_CDNS_719427747080 $T=56340 148580 0 0 $X=54830 $Y=147550
X1105 VDDA 6 6 pe3_CDNS_719427747080 $T=67580 148580 0 0 $X=66070 $Y=147550
X1106 VDDA 6 7 pe3_CDNS_719427747080 $T=78820 148580 0 0 $X=77310 $Y=147550
X1107 VDDA 6 6 pe3_CDNS_719427747080 $T=90060 148580 0 0 $X=88550 $Y=147550
X1108 VDDA 6 7 pe3_CDNS_719427747080 $T=101300 148580 0 0 $X=99790 $Y=147550
X1109 VDDA 6 6 pe3_CDNS_719427747080 $T=112540 148580 0 0 $X=111030 $Y=147550
X1110 VDDA 6 7 pe3_CDNS_719427747080 $T=123780 148580 0 0 $X=122270 $Y=147550
X1111 VDDA 6 6 pe3_CDNS_719427747080 $T=135020 148580 0 0 $X=133510 $Y=147550
X1112 VDDA 6 7 pe3_CDNS_719427747080 $T=146260 148580 0 0 $X=144750 $Y=147550
X1113 VDDA VDDA VDDA pe3_CDNS_719427747080 $T=157500 148580 0 0 $X=155990 $Y=147550
X1114 VDDA VDDA VDDA pe3_CDNS_719427747080 $T=362795 71115 1 0 $X=361285 $Y=60085
X1115 VDDA VDDA VDDA pe3_CDNS_719427747080 $T=362795 89915 1 0 $X=361285 $Y=78885
X1116 VDDA VDDA VDDA pe3_CDNS_719427747080 $T=362795 108715 1 0 $X=361285 $Y=97685
X1117 VDDA VDDA VDDA pe3_CDNS_719427747080 $T=362795 127515 1 0 $X=361285 $Y=116485
X1118 VDDA VDDA VDDA pe3_CDNS_719427747080 $T=362795 146315 1 0 $X=361285 $Y=135285
X1119 VDDA VDDA VDDA pe3_CDNS_719427747080 $T=362795 165115 1 0 $X=361285 $Y=154085
X1120 19 9 VOUT VDDA GNDA pe3_CDNS_719427747081 $T=373510 36320 1 0 $X=372000 $Y=25290
X1121 17 9 VOUT VDDA GNDA pe3_CDNS_719427747082 $T=364135 36320 1 0 $X=362625 $Y=25290
X1122 20 9 VOUT VDDA GNDA pe3_CDNS_719427747083 $T=351800 36320 1 0 $X=350290 $Y=25290
X1123 16 9 VOUT VDDA GNDA pe3_CDNS_719427747084 $T=333335 36320 1 0 $X=331825 $Y=25290
X1124 15 9 VOUT VDDA GNDA pe3_CDNS_719427747085 $T=302570 36320 1 0 $X=301060 $Y=25290
X1125 14 9 VOUT VDDA GNDA pe3_CDNS_719427747086 $T=246755 36320 1 0 $X=245245 $Y=25290
X1126 VOUT GNDA rpp1k1_3_CDNS_719427747087 $T=190390 9160 0 0 $X=185230 $Y=8940
X1127 18 9 21 VDDA GNDA pe3_CDNS_719427747088 $T=223935 36320 1 0 $X=222425 $Y=25290
X1128 21 GNDA rpp1k1_3_CDNS_719427747089 $T=80195 9200 0 0 $X=75035 $Y=8980
X1129 8 GNDA GNDA pe3_CDNS_7194277470810 $T=154675 76695 0 0 $X=153165 $Y=75665
X1130 9 8 GNDA pe3_CDNS_7194277470810 $T=154675 98175 0 0 $X=153165 $Y=97145
X1131 10 9 GNDA pe3_CDNS_7194277470810 $T=154675 119125 0 0 $X=153165 $Y=118095
X1132 VDDA ENABLE 31 pe3_CDNS_7194277470811 $T=91085 67915 1 0 $X=90175 $Y=61345
X1133 14 D5 GNDA VDDA pe3_CDNS_7194277470812 $T=307075 17335 1 0 $X=305565 $Y=6305
X1134 15 D4 GNDA VDDA pe3_CDNS_7194277470812 $T=316335 17335 1 0 $X=314825 $Y=6305
X1135 16 D3 GNDA VDDA pe3_CDNS_7194277470812 $T=325595 17335 1 0 $X=324085 $Y=6305
X1136 20 D2 GNDA VDDA pe3_CDNS_7194277470812 $T=334855 17335 1 0 $X=333345 $Y=6305
X1137 17 D1 GNDA VDDA pe3_CDNS_7194277470812 $T=344115 17335 1 0 $X=342605 $Y=6305
X1138 19 D0 GNDA VDDA pe3_CDNS_7194277470812 $T=353375 17335 1 0 $X=351865 $Y=6305
X1139 1 BIAS BIAS GNDA ne3_CDNS_7194277470813 $T=7715 59435 0 0 $X=6915 $Y=59035
X1140 3 BIAS 4 GNDA ne3_CDNS_7194277470813 $T=34470 59435 0 0 $X=33670 $Y=59035
X1141 12 BIAS 13 GNDA ne3_CDNS_7194277470813 $T=62205 59435 0 0 $X=61405 $Y=59035
X1142 GNDA GNDA GNDA ne3_CDNS_7194277470815 $T=11530 16320 0 0 $X=10730 $Y=15920
X1143 GNDA GNDA GNDA ne3_CDNS_7194277470815 $T=11530 38460 1 0 $X=10730 $Y=27890
X1144 GNDA 1 12 ne3_CDNS_7194277470815 $T=14770 16320 0 0 $X=13970 $Y=15920
X1145 GNDA 1 1 ne3_CDNS_7194277470815 $T=14770 38460 1 0 $X=13970 $Y=27890
X1146 GNDA 1 3 ne3_CDNS_7194277470815 $T=18010 16320 0 0 $X=17210 $Y=15920
X1147 GNDA 1 12 ne3_CDNS_7194277470815 $T=18010 38460 1 0 $X=17210 $Y=27890
X1148 GNDA 1 1 ne3_CDNS_7194277470815 $T=21250 16320 0 0 $X=20450 $Y=15920
X1149 GNDA 1 3 ne3_CDNS_7194277470815 $T=21250 38460 1 0 $X=20450 $Y=27890
X1150 GNDA 1 12 ne3_CDNS_7194277470815 $T=24490 16320 0 0 $X=23690 $Y=15920
X1151 GNDA 1 1 ne3_CDNS_7194277470815 $T=24490 38460 1 0 $X=23690 $Y=27890
X1152 GNDA 1 3 ne3_CDNS_7194277470815 $T=27730 16320 0 0 $X=26930 $Y=15920
X1153 GNDA 1 12 ne3_CDNS_7194277470815 $T=27730 38460 1 0 $X=26930 $Y=27890
X1154 GNDA 1 1 ne3_CDNS_7194277470815 $T=30970 16320 0 0 $X=30170 $Y=15920
X1155 GNDA 1 3 ne3_CDNS_7194277470815 $T=30970 38460 1 0 $X=30170 $Y=27890
X1156 GNDA 1 12 ne3_CDNS_7194277470815 $T=34210 16320 0 0 $X=33410 $Y=15920
X1157 GNDA 1 1 ne3_CDNS_7194277470815 $T=34210 38460 1 0 $X=33410 $Y=27890
X1158 GNDA 1 3 ne3_CDNS_7194277470815 $T=37450 16320 0 0 $X=36650 $Y=15920
X1159 GNDA 1 12 ne3_CDNS_7194277470815 $T=37450 38460 1 0 $X=36650 $Y=27890
X1160 GNDA 1 1 ne3_CDNS_7194277470815 $T=40690 16320 0 0 $X=39890 $Y=15920
X1161 GNDA 1 3 ne3_CDNS_7194277470815 $T=40690 38460 1 0 $X=39890 $Y=27890
X1162 GNDA 1 12 ne3_CDNS_7194277470815 $T=43930 16320 0 0 $X=43130 $Y=15920
X1163 GNDA 1 1 ne3_CDNS_7194277470815 $T=43930 38460 1 0 $X=43130 $Y=27890
X1164 GNDA 1 3 ne3_CDNS_7194277470815 $T=47170 16320 0 0 $X=46370 $Y=15920
X1165 GNDA 1 12 ne3_CDNS_7194277470815 $T=47170 38460 1 0 $X=46370 $Y=27890
X1166 GNDA 1 1 ne3_CDNS_7194277470815 $T=50410 16320 0 0 $X=49610 $Y=15920
X1167 GNDA 1 3 ne3_CDNS_7194277470815 $T=50410 38460 1 0 $X=49610 $Y=27890
X1168 GNDA GNDA GNDA ne3_CDNS_7194277470815 $T=53650 16320 0 0 $X=52850 $Y=15920
X1169 GNDA GNDA GNDA ne3_CDNS_7194277470815 $T=53650 38460 1 0 $X=52850 $Y=27890
X1170 VDDA pe3_CDNS_7194277470816 $T=362795 52315 1 0 $X=361285 $Y=49285
X1171 VDDA pe3_CDNS_7194277470816 $T=362795 175915 1 0 $X=361285 $Y=172885
X1172 GNDA 31 1 ne3_CDNS_7194277470817 $T=96785 56345 0 0 $X=95985 $Y=55765
X1173 GNDA 31 VOUT ne3_CDNS_7194277470817 $T=102390 56345 0 0 $X=101590 $Y=55765
X1174 GNDA ENABLE 31 ne3_CDNS_7194277470818 $T=91035 56560 0 0 $X=90235 $Y=56160
X1175 VDDA MASCO__A1 $T=203925 49285 0 0 $X=203925 $Y=49285
X1176 VDDA MASCO__A1 $T=203925 172885 0 0 $X=203925 $Y=172885
X1177 VDDA MASCO__A1 $T=226405 49285 0 0 $X=226405 $Y=49285
X1178 VDDA MASCO__A1 $T=226405 172885 0 0 $X=226405 $Y=172885
X1179 VDDA MASCO__A1 $T=248885 49285 0 0 $X=248885 $Y=49285
X1180 VDDA MASCO__A1 $T=248885 172885 0 0 $X=248885 $Y=172885
X1181 VDDA MASCO__A1 $T=271365 49285 0 0 $X=271365 $Y=49285
X1182 VDDA MASCO__A1 $T=271365 172885 0 0 $X=271365 $Y=172885
X1183 VDDA MASCO__A1 $T=293845 49285 0 0 $X=293845 $Y=49285
X1184 VDDA MASCO__A1 $T=293845 172885 0 0 $X=293845 $Y=172885
X1185 VDDA MASCO__A1 $T=316325 49285 0 0 $X=316325 $Y=49285
X1186 VDDA MASCO__A1 $T=316325 172885 0 0 $X=316325 $Y=172885
X1187 VDDA MASCO__A1 $T=338805 49285 0 0 $X=338805 $Y=49285
X1188 VDDA MASCO__A1 $T=338805 172885 0 0 $X=338805 $Y=172885
X1189 VDDA 10 4 4 4 MASCO__A2 $T=14200 160530 0 0 $X=14200 $Y=160530
X1190 VDDA 6 VDDA 6 VDDA MASCO__A2 $T=144750 160530 0 0 $X=144750 $Y=160530
X1191 VDDA VDDA VDDA VDDA VDDA MASCO__A2 $T=338805 60085 0 0 $X=338805 $Y=60085
X1192 VDDA 14 14 7 7 MASCO__A2 $T=338805 78885 0 0 $X=338805 $Y=78885
X1193 VDDA 14 14 7 7 MASCO__A2 $T=338805 97685 0 0 $X=338805 $Y=97685
X1194 VDDA 14 14 7 7 MASCO__A2 $T=338805 116485 0 0 $X=338805 $Y=116485
X1195 VDDA 14 14 7 7 MASCO__A2 $T=338805 135285 0 0 $X=338805 $Y=135285
X1196 VDDA 14 14 7 7 MASCO__A2 $T=338805 154085 0 0 $X=338805 $Y=154085
X1197 13 VDDA 13 13 7 6 21 13 VREF 13
+ GNDA MASCO__B5 $T=66310 96535 0 0 $X=66310 $Y=96535
X1198 13 VDDA 6 7 7 6 21 VREF VREF 21
+ GNDA MASCO__B5 $T=73110 96535 0 0 $X=73110 $Y=96535
X1199 13 VDDA 6 7 7 6 21 VREF VREF 21
+ GNDA MASCO__B5 $T=79910 96535 0 0 $X=79910 $Y=96535
X1200 13 VDDA 6 7 7 6 21 VREF VREF 21
+ GNDA MASCO__B5 $T=86710 96535 0 0 $X=86710 $Y=96535
X1201 13 VDDA 6 7 7 6 21 VREF VREF 21
+ GNDA MASCO__B5 $T=93510 96535 0 0 $X=93510 $Y=96535
X1202 13 VDDA 6 7 7 6 21 VREF VREF 21
+ GNDA MASCO__B5 $T=100310 96535 0 0 $X=100310 $Y=96535
X1203 13 VDDA 6 7 7 6 21 VREF VREF 21
+ GNDA MASCO__B5 $T=107110 96535 0 0 $X=107110 $Y=96535
X1204 13 VDDA 6 7 7 6 21 VREF VREF 21
+ GNDA MASCO__B5 $T=113910 96535 0 0 $X=113910 $Y=96535
X1205 13 VDDA 6 7 13 13 13 VREF 13 21
+ GNDA MASCO__B5 $T=120710 96535 0 0 $X=120710 $Y=96535
X1206 VDDA VDDA 6 7 6 7 VDDA MASCO__A6 $T=54830 160530 0 0 $X=54830 $Y=160530
X1207 VDDA 6 6 7 6 7 6 MASCO__A6 $T=99790 160530 0 0 $X=99790 $Y=160530
X1208 VDDA VDDA 7 14 15 15 VDDA MASCO__A6 $T=203925 60085 0 0 $X=203925 $Y=60085
X1209 VDDA VDDA 7 14 15 16 VDDA MASCO__A6 $T=203925 78885 0 0 $X=203925 $Y=78885
X1210 VDDA VDDA 7 14 15 16 VDDA MASCO__A6 $T=203925 97685 0 0 $X=203925 $Y=97685
X1211 VDDA VDDA 7 14 15 16 VDDA MASCO__A6 $T=203925 116485 0 0 $X=203925 $Y=116485
X1212 VDDA VDDA 7 14 15 16 VDDA MASCO__A6 $T=203925 135285 0 0 $X=203925 $Y=135285
X1213 VDDA VDDA 7 14 14 14 VDDA MASCO__A6 $T=203925 154085 0 0 $X=203925 $Y=154085
X1214 VDDA 15 7 15 18 14 7 MASCO__A6 $T=248885 60085 0 0 $X=248885 $Y=60085
X1215 VDDA 18 7 20 20 18 7 MASCO__A6 $T=248885 78885 0 0 $X=248885 $Y=78885
X1216 VDDA 17 7 18 19 18 7 MASCO__A6 $T=248885 97685 0 0 $X=248885 $Y=97685
X1217 VDDA 18 7 17 18 16 7 MASCO__A6 $T=248885 116485 0 0 $X=248885 $Y=116485
X1218 VDDA 18 7 20 20 18 7 MASCO__A6 $T=248885 135285 0 0 $X=248885 $Y=135285
X1219 VDDA 14 7 14 15 15 7 MASCO__A6 $T=248885 154085 0 0 $X=248885 $Y=154085
X1220 VDDA 14 VDDA VDDA VDDA VDDA 7 MASCO__A6 $T=293845 60085 0 0 $X=293845 $Y=60085
X1221 VDDA 16 7 15 14 14 7 MASCO__A6 $T=293845 78885 0 0 $X=293845 $Y=78885
X1222 VDDA 16 7 15 14 14 7 MASCO__A6 $T=293845 97685 0 0 $X=293845 $Y=97685
X1223 VDDA 15 7 15 14 14 7 MASCO__A6 $T=293845 116485 0 0 $X=293845 $Y=116485
X1224 VDDA 16 7 15 14 14 7 MASCO__A6 $T=293845 135285 0 0 $X=293845 $Y=135285
X1225 VDDA 15 7 18 14 14 7 MASCO__A6 $T=293845 154085 0 0 $X=293845 $Y=154085
D0 GNDA VDDA p_dnw AREA=7.95604e-10 PJ=0.00014876 perimeter=0.00014876 $X=8500 $Y=140710 $dt=3
D1 GNDA VDDA p_dnw AREA=2.14716e-09 PJ=0.0003306 perimeter=0.0003306 $X=48630 $Y=140710 $dt=3
D2 GNDA VDDA p_dnw AREA=3.11448e-11 PJ=3.188e-05 perimeter=3.188e-05 $X=88435 $Y=59745 $dt=3
D3 GNDA 8 p_dnw AREA=1.97548e-10 PJ=8.944e-05 perimeter=8.944e-05 $X=151005 $Y=72505 $dt=3
D4 GNDA 9 p_dnw AREA=1.97548e-10 PJ=8.944e-05 perimeter=8.944e-05 $X=151005 $Y=93985 $dt=3
D5 GNDA 10 p_dnw AREA=1.97548e-10 PJ=8.944e-05 perimeter=8.944e-05 $X=151005 $Y=114935 $dt=3
D6 GNDA VDDA p_dnw AREA=1.47356e-08 PJ=0.0006944 perimeter=0.0006944 $X=181765 $Y=46865 $dt=3
D7 GNDA VDDA p_dnw AREA=1.65707e-09 PJ=0.00035483 perimeter=0.00035483 $X=220785 $Y=22870 $dt=3
D8 GNDA VDDA p_dnw AREA=6.02548e-10 PJ=0.00014223 perimeter=0.00014223 $X=303405 $Y=4665 $dt=3
D9 GNDA VDDA p_ddnw AREA=1.72778e-09 PJ=0.0002104 perimeter=0.0002104 $X=65040 $Y=95265 $dt=4
D10 13 VDDA p_dipdnwmv AREA=9.7703e-10 PJ=0.0001796 perimeter=0.0001796 $X=68890 $Y=99115 $dt=5
D11 GNDA VDDA p_dnw3 AREA=2.92576e-10 PJ=0 perimeter=0 $X=14200 $Y=147550 $dt=6
D12 GNDA VDDA p_dnw3 AREA=2.92576e-10 PJ=0 perimeter=0 $X=14200 $Y=160530 $dt=6
D13 GNDA VDDA p_dnw3 AREA=1.37701e-09 PJ=0 perimeter=0 $X=54830 $Y=147550 $dt=6
D14 GNDA VDDA p_dnw3 AREA=1.37701e-09 PJ=0 perimeter=0 $X=54830 $Y=160530 $dt=6
D15 GNDA VDDA p_dnw3 AREA=2.67592e-11 PJ=0 perimeter=0 $X=89575 $Y=60885 $dt=6
D16 GNDA VDDA p_dnw3 AREA=6.91743e-10 PJ=0 perimeter=0 $X=203925 $Y=49285 $dt=6
D17 GNDA VDDA p_dnw3 AREA=2.05478e-09 PJ=0 perimeter=0 $X=203925 $Y=60085 $dt=6
D18 GNDA VDDA p_dnw3 AREA=2.05478e-09 PJ=0 perimeter=0 $X=203925 $Y=78885 $dt=6
D19 GNDA VDDA p_dnw3 AREA=2.05478e-09 PJ=0 perimeter=0 $X=203925 $Y=97685 $dt=6
D20 GNDA VDDA p_dnw3 AREA=2.05478e-09 PJ=0 perimeter=0 $X=203925 $Y=116485 $dt=6
D21 GNDA VDDA p_dnw3 AREA=2.05478e-09 PJ=0 perimeter=0 $X=203925 $Y=135285 $dt=6
D22 GNDA VDDA p_dnw3 AREA=2.05478e-09 PJ=0 perimeter=0 $X=203925 $Y=154085 $dt=6
D23 GNDA VDDA p_dnw3 AREA=6.91743e-10 PJ=0 perimeter=0 $X=203925 $Y=172885 $dt=6
.ends dac6b_amp_n2
