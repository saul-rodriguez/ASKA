* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : current_source_gm_10_en_r                    *
* Netlisted  : Tue Aug 13 03:37:13 2024                     *
* PVS Version: 23.10-p043 Mon Oct 2 18:09:08 PDT 2023      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 LDDN(nedia) nedia2_d dnwtrm(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 1 MN(ne3) nem ndiff(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 2 MP(pe3) pem pdiff(D) p1trm(G) pdiff(S) nwtrm(B)
*.DEVTMPLT 3 MOSVC3() mosvcm p1trm(G) nwtrm(NW) bulk(SB)
*.DEVTMPLT 4 R(s_res) s_res bulk(POS) bulk(NEG)
*.DEVTMPLT 5 D(p_dnw) p_dnw bulk(POS) nwtrm(NEG)
*.DEVTMPLT 6 D(p_dnw3) p_dnwm bulk(POS) nwtrm(NEG)
*.DEVTMPLT 7 R(rpp1k1_3) rpp1k1_s p1trm(POS) p1trm(NEG) bulk(SUB)
*.DEVTMPLT 8 R(rpp1k1_3) rpp1k1_n p1trm(POS) p1trm(NEG) nwtrm(SUB)
*.DEVTMPLT 9 C(cmm5t) cmim capm(POS) m4trm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MOSVC3                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MOSVC3 G NW SB
.ends MOSVC3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: LDDN                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt LDDN D G S B
.ends LDDN

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_723534627840                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_723534627840 1 2 3
** N=3 EP=3 FDC=4
M0 3 2 1 1 ne3 L=5e-07 W=5e-06 AD=1.35e-12 AS=2.4e-12 PD=5.54e-06 PS=1.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 1 ne3 L=5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=1040 $Y=0 $dt=1
M2 3 2 1 1 ne3 L=5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=2080 $Y=0 $dt=1
M3 1 2 3 1 ne3 L=5e-07 W=5e-06 AD=2.4e-12 AS=1.35e-12 PD=1.096e-05 PS=5.54e-06 $X=3120 $Y=0 $dt=1
.ends ne3_CDNS_723534627840

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nedia_CDNS_723534627841                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nedia_CDNS_723534627841 1 2 3 4
** N=4 EP=4 FDC=1
X0 2 4 3 1 LDDN w=5e-05 l=1.25e-06 adio=1.08602e-09 pdio=0.00013535 extlay=1 $[nedia] $X=-680 $Y=-4850 $dt=0
.ends nedia_CDNS_723534627841

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_723534627842                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_723534627842 1 2 3
** N=3 EP=3 FDC=4
M0 3 2 1 1 ne3 L=3.5e-07 W=5e-06 AD=1.35e-12 AS=2.4e-12 PD=5.54e-06 PS=1.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 1 ne3 L=3.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=890 $Y=0 $dt=1
M2 3 2 1 1 ne3 L=3.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=1780 $Y=0 $dt=1
M3 1 2 3 1 ne3 L=3.5e-07 W=5e-06 AD=2.4e-12 AS=1.35e-12 PD=1.096e-05 PS=5.54e-06 $X=2670 $Y=0 $dt=1
.ends ne3_CDNS_723534627842

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_723534627843                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_723534627843 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.00010265 W=4e-06 $[rpp1k1_3] $SUB=3 $X=0 $Y=0 $dt=7
.ends rpp1k1_3_CDNS_723534627843

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nedia_CDNS_723534627844                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nedia_CDNS_723534627844 1 2 3 4
** N=4 EP=4 FDC=8
X0 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=-680 $Y=-4850 $dt=0
X1 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=11220 $Y=-4850 $dt=0
X2 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=23120 $Y=-4850 $dt=0
X3 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=35020 $Y=-4850 $dt=0
X4 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=46920 $Y=-4850 $dt=0
X5 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=58820 $Y=-4850 $dt=0
X6 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=70720 $Y=-4850 $dt=0
X7 2 4 3 1 LDDN w=0.0001 l=1.25e-06 adio=1.01941e-09 pdio=4.39938e-05 extlay=1 $[nedia] $X=82620 $Y=-4850 $dt=0
.ends nedia_CDNS_723534627844

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_723534627845                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_723534627845 1 2 3 4
** N=4 EP=4 FDC=2
M0 3 2 1 4 ne3 L=1e-05 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 ne3 L=1e-05 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=10540 $Y=0 $dt=1
.ends ne3_CDNS_723534627845

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_723534627846                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_723534627846 1 2 3
*.DEVICECLIMB
** N=4 EP=3 FDC=1
M0 3 2 1 1 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
.ends pe3_CDNS_723534627846

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_723534627847                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_723534627847 1 2 3
*.DEVICECLIMB
** N=4 EP=3 FDC=2
M0 3 2 1 1 pe3 L=3e-07 W=3e-06 AD=8.1e-13 AS=1.44e-12 PD=3.54e-06 PS=6.96e-06 $X=0 $Y=0 $dt=2
M1 1 2 3 1 pe3 L=3e-07 W=3e-06 AD=1.44e-12 AS=8.1e-13 PD=6.96e-06 PS=3.54e-06 $X=840 $Y=0 $dt=2
.ends pe3_CDNS_723534627847

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_723534627848                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_723534627848 1 2 3
** N=3 EP=3 FDC=1
R0 1 2 L=0.00204354 W=2e-06 $[rpp1k1_3] $SUB=3 $X=-2220 $Y=0 $dt=7
.ends rpp1k1_3_CDNS_723534627848

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7235346278411                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7235346278411 1 2 3 4
*.DEVICECLIMB
** N=5 EP=4 FDC=1
M0 3 2 1 4 pe3 L=5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
.ends pe3_CDNS_7235346278411

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7235346278412                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7235346278412 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=1e-05 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends ne3_CDNS_7235346278412

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7235346278413                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7235346278413 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=1e-06 W=5e-06 AD=2.4e-12 AS=2.4e-12 PD=1.096e-05 PS=1.096e-05 $X=0 $Y=0 $dt=1
.ends ne3_CDNS_7235346278413

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7235346278414                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7235346278414 1 2 3
*.DEVICECLIMB
** N=3 EP=3 FDC=9
M0 3 2 1 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=2
M1 1 2 3 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=5540 $Y=0 $dt=2
M2 3 2 1 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=11080 $Y=0 $dt=2
M3 1 2 3 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=16620 $Y=0 $dt=2
M4 3 2 1 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=22160 $Y=0 $dt=2
M5 1 2 3 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=27700 $Y=0 $dt=2
M6 3 2 1 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=33240 $Y=0 $dt=2
M7 1 2 3 1 pe3 L=5e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=38780 $Y=0 $dt=2
M8 3 2 1 1 pe3 L=5e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=44320 $Y=0 $dt=2
.ends pe3_CDNS_7235346278414

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7235346278415                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7235346278415 1 2 3
** N=3 EP=3 FDC=1
R0 1 2 L=1e-05 W=2e-06 $[rpp1k1_3] $SUB=3 $X=0 $Y=0 $dt=7
.ends rpp1k1_3_CDNS_7235346278415

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7235346278416                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7235346278416 1 2 3
*.DEVICECLIMB
** N=4 EP=3 FDC=1
R0 2 1 L=0.00016435 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=8
.ends rpp1k1_3_CDNS_7235346278416

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7235346278417                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7235346278417 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.00041122 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=7
.ends rpp1k1_3_CDNS_7235346278417

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7235346278418                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7235346278418 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=3.5e-07 W=2e-06 AD=9.6e-13 AS=9.6e-13 PD=4.96e-06 PS=4.96e-06 $X=0 $Y=0 $dt=1
.ends ne3_CDNS_7235346278418

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: current_source_gm_10_en_r                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt current_source_gm_10_en_r BIAS EN FB GNDA GNDHV IN OUT PACTIVE VDD3A VDDHV
+ VSUBHV
** N=27 EP=11 FDC=198
X399 GNDA 11 10 ne3_CDNS_723534627840 $T=248120 21400 0 0 $X=247320 $Y=21000
X400 VSUBHV 15 GNDHV 10 nedia_CDNS_723534627841 $T=282450 37820 0 0 $X=266230 $Y=18430
X401 GNDA 22 1 ne3_CDNS_723534627842 $T=25060 81535 0 0 $X=24260 $Y=80955
X402 GNDA 21 11 ne3_CDNS_723534627842 $T=30635 81535 0 0 $X=29835 $Y=80955
X403 15 GNDHV VSUBHV rpp1k1_3_CDNS_723534627843 $T=317545 27490 0 90 $X=309065 $Y=26550
X404 VSUBHV OUT FB 15 nedia_CDNS_723534627844 $T=441980 141045 0 270 $X=422590 $Y=41525
X405 1 BIAS BIAS GNDA ne3_CDNS_723534627845 $T=8060 64240 0 0 $X=7260 $Y=63840
X406 3 BIAS 4 GNDA ne3_CDNS_723534627845 $T=33845 64240 0 0 $X=33045 $Y=63840
X407 5 BIAS 6 GNDA ne3_CDNS_723534627845 $T=59570 64240 0 0 $X=58770 $Y=63840
X408 VDD3A 4 10 pe3_CDNS_723534627846 $T=63965 94930 0 180 $X=61455 $Y=83900
X409 VDD3A 4 10 pe3_CDNS_723534627846 $T=66205 94930 0 180 $X=63695 $Y=83900
X410 VDD3A 4 4 pe3_CDNS_723534627846 $T=68445 94930 0 180 $X=65935 $Y=83900
X411 VDD3A 4 10 pe3_CDNS_723534627846 $T=70685 94930 0 180 $X=68175 $Y=83900
X412 VDD3A 4 10 pe3_CDNS_723534627846 $T=72925 94930 0 180 $X=70415 $Y=83900
X413 VDD3A EN 22 pe3_CDNS_723534627847 $T=15530 89865 0 180 $X=13480 $Y=86295
X414 VDD3A PACTIVE 21 pe3_CDNS_723534627847 $T=19690 89865 0 180 $X=17640 $Y=86295
X415 GNDHV OUT VSUBHV rpp1k1_3_CDNS_723534627848 $T=558265 45130 0 90 $X=515365 $Y=41970
X416 VDD3A VDD3A VDD3A VDD3A pe3_CDNS_7235346278411 $T=109700 69700 0 0 $X=108190 $Y=68670
X417 VDD3A VDD3A VDD3A VDD3A pe3_CDNS_7235346278411 $T=109700 93320 1 0 $X=108190 $Y=82290
X418 VDD3A VDD3A VDD3A VDD3A pe3_CDNS_7235346278411 $T=113660 125985 0 0 $X=112150 $Y=124955
X419 VDD3A VDD3A VDD3A VDD3A pe3_CDNS_7235346278411 $T=113660 148965 1 0 $X=112150 $Y=137935
X420 13 8 11 VDD3A pe3_CDNS_7235346278411 $T=115940 69700 0 0 $X=114430 $Y=68670
X421 13 7 12 VDD3A pe3_CDNS_7235346278411 $T=115940 93320 1 0 $X=114430 $Y=82290
X422 VDD3A 6 13 VDD3A pe3_CDNS_7235346278411 $T=119900 125985 0 0 $X=118390 $Y=124955
X423 VDD3A 6 13 VDD3A pe3_CDNS_7235346278411 $T=119900 148965 1 0 $X=118390 $Y=137935
X424 13 7 12 VDD3A pe3_CDNS_7235346278411 $T=122180 69700 0 0 $X=120670 $Y=68670
X425 13 8 11 VDD3A pe3_CDNS_7235346278411 $T=122180 93320 1 0 $X=120670 $Y=82290
X426 VDD3A 6 13 VDD3A pe3_CDNS_7235346278411 $T=126140 125985 0 0 $X=124630 $Y=124955
X427 VDD3A 6 13 VDD3A pe3_CDNS_7235346278411 $T=126140 148965 1 0 $X=124630 $Y=137935
X428 13 8 11 VDD3A pe3_CDNS_7235346278411 $T=128420 69700 0 0 $X=126910 $Y=68670
X429 13 7 12 VDD3A pe3_CDNS_7235346278411 $T=128420 93320 1 0 $X=126910 $Y=82290
X430 VDD3A 6 13 VDD3A pe3_CDNS_7235346278411 $T=132380 125985 0 0 $X=130870 $Y=124955
X431 VDD3A 6 13 VDD3A pe3_CDNS_7235346278411 $T=132380 148965 1 0 $X=130870 $Y=137935
X432 13 7 12 VDD3A pe3_CDNS_7235346278411 $T=134660 69700 0 0 $X=133150 $Y=68670
X433 13 8 11 VDD3A pe3_CDNS_7235346278411 $T=134660 93320 1 0 $X=133150 $Y=82290
X434 VDD3A 6 13 VDD3A pe3_CDNS_7235346278411 $T=138620 125985 0 0 $X=137110 $Y=124955
X435 VDD3A 6 13 VDD3A pe3_CDNS_7235346278411 $T=138620 148965 1 0 $X=137110 $Y=137935
X436 13 8 11 VDD3A pe3_CDNS_7235346278411 $T=140900 69700 0 0 $X=139390 $Y=68670
X437 13 7 12 VDD3A pe3_CDNS_7235346278411 $T=140900 93320 1 0 $X=139390 $Y=82290
X438 VDD3A 6 13 VDD3A pe3_CDNS_7235346278411 $T=144860 125985 0 0 $X=143350 $Y=124955
X439 VDD3A 6 13 VDD3A pe3_CDNS_7235346278411 $T=144860 148965 1 0 $X=143350 $Y=137935
X440 13 7 12 VDD3A pe3_CDNS_7235346278411 $T=147140 69700 0 0 $X=145630 $Y=68670
X441 13 8 11 VDD3A pe3_CDNS_7235346278411 $T=147140 93320 1 0 $X=145630 $Y=82290
X442 VDD3A 6 8 VDD3A pe3_CDNS_7235346278411 $T=151100 125985 0 0 $X=149590 $Y=124955
X443 VDD3A 6 7 VDD3A pe3_CDNS_7235346278411 $T=151100 148965 1 0 $X=149590 $Y=137935
X444 13 8 11 VDD3A pe3_CDNS_7235346278411 $T=153380 69700 0 0 $X=151870 $Y=68670
X445 13 7 12 VDD3A pe3_CDNS_7235346278411 $T=153380 93320 1 0 $X=151870 $Y=82290
X446 VDD3A 6 6 VDD3A pe3_CDNS_7235346278411 $T=157340 125985 0 0 $X=155830 $Y=124955
X447 VDD3A 6 6 VDD3A pe3_CDNS_7235346278411 $T=157340 148965 1 0 $X=155830 $Y=137935
X448 13 7 12 VDD3A pe3_CDNS_7235346278411 $T=159620 69700 0 0 $X=158110 $Y=68670
X449 13 8 11 VDD3A pe3_CDNS_7235346278411 $T=159620 93320 1 0 $X=158110 $Y=82290
X450 VDD3A 6 7 VDD3A pe3_CDNS_7235346278411 $T=163580 125985 0 0 $X=162070 $Y=124955
X451 VDD3A 6 8 VDD3A pe3_CDNS_7235346278411 $T=163580 148965 1 0 $X=162070 $Y=137935
X452 13 8 11 VDD3A pe3_CDNS_7235346278411 $T=165860 69700 0 0 $X=164350 $Y=68670
X453 13 7 12 VDD3A pe3_CDNS_7235346278411 $T=165860 93320 1 0 $X=164350 $Y=82290
X454 VDD3A 6 13 VDD3A pe3_CDNS_7235346278411 $T=169820 125985 0 0 $X=168310 $Y=124955
X455 VDD3A 6 13 VDD3A pe3_CDNS_7235346278411 $T=169820 148965 1 0 $X=168310 $Y=137935
X456 13 7 12 VDD3A pe3_CDNS_7235346278411 $T=172100 69700 0 0 $X=170590 $Y=68670
X457 13 8 11 VDD3A pe3_CDNS_7235346278411 $T=172100 93320 1 0 $X=170590 $Y=82290
X458 VDD3A 6 13 VDD3A pe3_CDNS_7235346278411 $T=176060 125985 0 0 $X=174550 $Y=124955
X459 VDD3A 6 13 VDD3A pe3_CDNS_7235346278411 $T=176060 148965 1 0 $X=174550 $Y=137935
X460 13 8 11 VDD3A pe3_CDNS_7235346278411 $T=178340 69700 0 0 $X=176830 $Y=68670
X461 13 7 12 VDD3A pe3_CDNS_7235346278411 $T=178340 93320 1 0 $X=176830 $Y=82290
X462 VDD3A 6 13 VDD3A pe3_CDNS_7235346278411 $T=182300 125985 0 0 $X=180790 $Y=124955
X463 VDD3A 6 13 VDD3A pe3_CDNS_7235346278411 $T=182300 148965 1 0 $X=180790 $Y=137935
X464 13 7 12 VDD3A pe3_CDNS_7235346278411 $T=184580 69700 0 0 $X=183070 $Y=68670
X465 13 8 11 VDD3A pe3_CDNS_7235346278411 $T=184580 93320 1 0 $X=183070 $Y=82290
X466 VDD3A 6 13 VDD3A pe3_CDNS_7235346278411 $T=188540 125985 0 0 $X=187030 $Y=124955
X467 VDD3A 6 13 VDD3A pe3_CDNS_7235346278411 $T=188540 148965 1 0 $X=187030 $Y=137935
X468 13 8 11 VDD3A pe3_CDNS_7235346278411 $T=190820 69700 0 0 $X=189310 $Y=68670
X469 13 7 12 VDD3A pe3_CDNS_7235346278411 $T=190820 93320 1 0 $X=189310 $Y=82290
X470 VDD3A 6 13 VDD3A pe3_CDNS_7235346278411 $T=194780 125985 0 0 $X=193270 $Y=124955
X471 VDD3A 6 13 VDD3A pe3_CDNS_7235346278411 $T=194780 148965 1 0 $X=193270 $Y=137935
X472 13 7 12 VDD3A pe3_CDNS_7235346278411 $T=197060 69700 0 0 $X=195550 $Y=68670
X473 13 8 11 VDD3A pe3_CDNS_7235346278411 $T=197060 93320 1 0 $X=195550 $Y=82290
X474 VDD3A VDD3A VDD3A VDD3A pe3_CDNS_7235346278411 $T=201020 125985 0 0 $X=199510 $Y=124955
X475 VDD3A VDD3A VDD3A VDD3A pe3_CDNS_7235346278411 $T=201020 148965 1 0 $X=199510 $Y=137935
X476 VDD3A VDD3A VDD3A VDD3A pe3_CDNS_7235346278411 $T=203300 69700 0 0 $X=201790 $Y=68670
X477 VDD3A VDD3A VDD3A VDD3A pe3_CDNS_7235346278411 $T=203300 93320 1 0 $X=201790 $Y=82290
X478 GNDA GNDA GNDA ne3_CDNS_7235346278412 $T=17420 20740 0 0 $X=16620 $Y=20340
X479 GNDA GNDA GNDA ne3_CDNS_7235346278412 $T=17420 42860 1 0 $X=16620 $Y=32290
X480 GNDA 1 5 ne3_CDNS_7235346278412 $T=28660 20740 0 0 $X=27860 $Y=20340
X481 GNDA 1 5 ne3_CDNS_7235346278412 $T=28660 42860 1 0 $X=27860 $Y=32290
X482 GNDA 1 1 ne3_CDNS_7235346278412 $T=39900 20740 0 0 $X=39100 $Y=20340
X483 GNDA 1 1 ne3_CDNS_7235346278412 $T=39900 42860 1 0 $X=39100 $Y=32290
X484 GNDA 1 3 ne3_CDNS_7235346278412 $T=51140 20740 0 0 $X=50340 $Y=20340
X485 GNDA 1 3 ne3_CDNS_7235346278412 $T=51140 42860 1 0 $X=50340 $Y=32290
X486 GNDA GNDA GNDA ne3_CDNS_7235346278412 $T=62380 20740 0 0 $X=61580 $Y=20340
X487 GNDA GNDA GNDA ne3_CDNS_7235346278412 $T=62380 42860 1 0 $X=61580 $Y=32290
X488 GNDA 12 11 ne3_CDNS_7235346278413 $T=232175 21040 0 0 $X=231375 $Y=20640
X489 GNDA 12 12 ne3_CDNS_7235346278413 $T=232175 32430 1 0 $X=231375 $Y=26860
X490 GNDA 12 12 ne3_CDNS_7235346278413 $T=234415 21040 0 0 $X=233615 $Y=20640
X491 GNDA 12 11 ne3_CDNS_7235346278413 $T=234415 32430 1 0 $X=233615 $Y=26860
X492 7 IN GNDA pe3_CDNS_7235346278414 $T=106815 19890 0 0 $X=105305 $Y=18860
X493 8 17 GNDA pe3_CDNS_7235346278414 $T=106815 43890 1 0 $X=105305 $Y=32860
X494 8 17 GNDA pe3_CDNS_7235346278414 $T=161095 19890 0 0 $X=159585 $Y=18860
X495 7 IN GNDA pe3_CDNS_7235346278414 $T=161095 43890 1 0 $X=159585 $Y=32860
X496 FB 17 GNDA rpp1k1_3_CDNS_7235346278415 $T=229190 61300 0 90 $X=226970 $Y=60360
X497 FB 17 GNDA rpp1k1_3_CDNS_7235346278415 $T=232060 61300 0 90 $X=229840 $Y=60360
X498 FB 17 GNDA rpp1k1_3_CDNS_7235346278415 $T=234930 61300 0 90 $X=232710 $Y=60360
X499 FB 17 GNDA rpp1k1_3_CDNS_7235346278415 $T=237800 61300 0 90 $X=235580 $Y=60360
X500 FB 17 GNDA rpp1k1_3_CDNS_7235346278415 $T=240670 61300 0 90 $X=238450 $Y=60360
X501 FB 17 GNDA rpp1k1_3_CDNS_7235346278415 $T=243540 61300 0 90 $X=241320 $Y=60360
X502 FB 17 GNDA rpp1k1_3_CDNS_7235346278415 $T=246410 61300 0 90 $X=244190 $Y=60360
X503 FB 17 GNDA rpp1k1_3_CDNS_7235346278415 $T=249280 61300 0 90 $X=247060 $Y=60360
X504 FB 17 GNDA rpp1k1_3_CDNS_7235346278415 $T=252150 61300 0 90 $X=249930 $Y=60360
X505 10 26 VDD3A rpp1k1_3_CDNS_7235346278416 $T=255085 124550 0 180 $X=228430 $Y=99030
X506 VDDHV 15 VSUBHV rpp1k1_3_CDNS_7235346278417 $T=322885 76685 0 270 $X=322665 $Y=25845
X507 GNDA EN 22 ne3_CDNS_7235346278418 $T=14340 81020 0 0 $X=13540 $Y=80620
X508 GNDA PACTIVE 21 ne3_CDNS_7235346278418 $T=18500 81020 0 0 $X=17700 $Y=80620
X751 VDD3A GNDA GNDA MOSVC3 w=2e-05 l=3e-05 $X=16180 $Y=110530 $dt=3
X752 VDD3A GNDA GNDA MOSVC3 w=2e-05 l=3e-05 $X=16180 $Y=132530 $dt=3
X753 VDD3A GNDA GNDA MOSVC3 w=2e-05 l=3e-05 $X=48780 $Y=110530 $dt=3
X754 VDD3A GNDA GNDA MOSVC3 w=2e-05 l=3e-05 $X=48780 $Y=132530 $dt=3
R4 GNDA VSUBHV 5 $[s_res] $X=263280 $Y=3815 $dt=4
D5 GNDA VDD3A p_dnw AREA=3.57048e-11 PJ=3.588e-05 perimeter=3.588e-05 $X=11740 $Y=84695 $dt=5
D6 GNDA VDD3A p_dnw AREA=1.90124e-10 PJ=7.516e-05 perimeter=7.516e-05 $X=59815 $Y=81480 $dt=5
D7 GNDA VDD3A p_dnw AREA=1.58288e-09 PJ=0.00049318 perimeter=0.00049318 $X=99710 $Y=59910 $dt=5
D8 GNDA VDD3A p_dnw AREA=3.09086e-09 PJ=0.00032604 perimeter=0.00032604 $X=101390 $Y=114415 $dt=5
D9 GNDA 7 p_dnw AREA=1.82058e-10 PJ=5.826e-05 perimeter=5.826e-05 $X=105905 $Y=15300 $dt=5
D10 GNDA 8 p_dnw AREA=1.82058e-10 PJ=5.826e-05 perimeter=5.826e-05 $X=105905 $Y=44920 $dt=5
D11 GNDA 8 p_dnw AREA=1.82058e-10 PJ=5.826e-05 perimeter=5.826e-05 $X=160185 $Y=15300 $dt=5
D12 GNDA 7 p_dnw AREA=1.82058e-10 PJ=5.826e-05 perimeter=5.826e-05 $X=160185 $Y=44920 $dt=5
D13 GNDA VDD3A p_dnw AREA=8.36476e-09 PJ=0.0003905 perimeter=0.0003905 $X=226790 $Y=95600 $dt=5
D14 GNDA VDD3A p_dnw3 AREA=4.20992e-11 PJ=0 perimeter=0 $X=12880 $Y=85835 $dt=6
D15 GNDA GNDA p_dnw3 AREA=5.9176e-11 PJ=0.00010492 perimeter=0.00010492 $X=15380 $Y=110100 $dt=6
D16 GNDA GNDA p_dnw3 AREA=5.9176e-11 PJ=0.00010492 perimeter=0.00010492 $X=15380 $Y=132100 $dt=6
D17 GNDA GNDA p_dnw3 AREA=5.9176e-11 PJ=0.00010492 perimeter=0.00010492 $X=47980 $Y=110100 $dt=6
D18 GNDA GNDA p_dnw3 AREA=5.9176e-11 PJ=0.00010492 perimeter=0.00010492 $X=47980 $Y=132100 $dt=6
D19 GNDA VDD3A p_dnw3 AREA=1.56539e-10 PJ=0 perimeter=0 $X=61455 $Y=83900 $dt=6
D20 GNDA 7 p_dnw3 AREA=5.86064e-10 PJ=7.406e-05 perimeter=7.406e-05 $X=105905 $Y=18860 $dt=6
D21 GNDA 8 p_dnw3 AREA=5.86064e-10 PJ=7.406e-05 perimeter=7.406e-05 $X=105905 $Y=33460 $dt=6
D22 GNDA VDD3A p_dnw3 AREA=1.22554e-09 PJ=0 perimeter=0 $X=108190 $Y=68670 $dt=6
D23 GNDA VDD3A p_dnw3 AREA=1.15225e-09 PJ=0.00012214 perimeter=0.00012214 $X=108190 $Y=82290 $dt=6
D24 GNDA VDD3A p_dnw3 AREA=1.15028e-09 PJ=0 perimeter=0 $X=112150 $Y=124955 $dt=6
D25 GNDA VDD3A p_dnw3 AREA=1.15028e-09 PJ=0 perimeter=0 $X=112150 $Y=137935 $dt=6
D26 GNDA 8 p_dnw3 AREA=5.86064e-10 PJ=7.406e-05 perimeter=7.406e-05 $X=160185 $Y=18860 $dt=6
D27 GNDA 7 p_dnw3 AREA=5.86064e-10 PJ=7.406e-05 perimeter=7.406e-05 $X=160185 $Y=33460 $dt=6
C28 11 26 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=231620 $Y=128940 $dt=9
C29 11 26 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=263220 $Y=97740 $dt=9
C30 11 26 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=263220 $Y=128940 $dt=9
C31 11 26 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=294820 $Y=97740 $dt=9
C32 11 26 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=294820 $Y=128940 $dt=9
C33 11 26 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=326420 $Y=97740 $dt=9
C34 11 26 area=8.4e-10 perimeter=0.000116 $[cmm5t] $X=326420 $Y=128940 $dt=9
.ends current_source_gm_10_en_r
