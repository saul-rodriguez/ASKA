* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : hvswitch5                                    *
* Netlisted  : Wed Aug  7 16:31:02 2024                     *
* PVS Version: 23.10-p043 Mon Oct 2 18:09:08 PDT 2023      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 LDDN(nedia) nedia2_d dnwtrm(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 1 LDDP(ped) ped12_d pwitrm(D) p1trm(G) pdiff(S) bulk(B)
*.DEVTMPLT 2 MN(ne3) nem ndiff(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 3 MP(pe3) pem pdiff(D) p1trm(G) pdiff(S) nwtrm(B)
*.DEVTMPLT 4 D(p_dnw) p_dnw bulk(POS) nwtrm(NEG)
*.DEVTMPLT 5 D(p_ddnw) p_ddnw bulk(POS) dnwtrm(NEG)
*.DEVTMPLT 6 D(p_dwhn) p_dwhn bulk(POS) hnw(NEG)
*.DEVTMPLT 7 D(dpp20) dpp20 pwitrm(POS) dnwtrm(NEG)
*.DEVTMPLT 8 D(dsba) d_dsba d_dsdf(POS) hnw(NEG) bulk(SUB)
*.DEVTMPLT 9 D(p_dnw3) p_dnwm bulk(POS) nwtrm(NEG)
*.DEVTMPLT 10 R(rpp1k1_3) rpp1k1_s p1trm(POS) p1trm(NEG) bulk(SUB)
*.DEVTMPLT 11 C(csf4a) d_csf4a m1atrm(POS) m1btrm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7230626554116                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7230626554116 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7230626554116

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7230626554136                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7230626554136 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7230626554136

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7230626554137                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7230626554137 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7230626554137

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7230626554145                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7230626554145 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7230626554145

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7230626554149                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7230626554149 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7230626554149

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7230626554150                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7230626554150 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7230626554150

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7230626554151                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7230626554151 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7230626554151

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7230626554153                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7230626554153 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7230626554153

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7230626554154                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7230626554154 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7230626554154

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7230626554157                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7230626554157 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7230626554157

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7230626554158                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7230626554158 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7230626554158

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nedia_CDNS_723062655410                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nedia_CDNS_723062655410 1 2 3 4
** N=4 EP=4 FDC=12
X0 2 3 4 1 LDDN w=5e-05 l=1.25e-06 adio=6.71697e-10 pdio=3.30958e-05 extlay=1 $[nedia] $X=-680 $Y=-4850 $dt=0
X1 2 3 4 1 LDDN w=5e-05 l=1.25e-06 adio=6.71697e-10 pdio=3.30958e-05 extlay=1 $[nedia] $X=11220 $Y=-4850 $dt=0
X2 2 3 4 1 LDDN w=5e-05 l=1.25e-06 adio=6.71697e-10 pdio=3.30958e-05 extlay=1 $[nedia] $X=23120 $Y=-4850 $dt=0
X3 2 3 4 1 LDDN w=5e-05 l=1.25e-06 adio=6.71697e-10 pdio=3.30958e-05 extlay=1 $[nedia] $X=35020 $Y=-4850 $dt=0
X4 2 3 4 1 LDDN w=5e-05 l=1.25e-06 adio=6.71697e-10 pdio=3.30958e-05 extlay=1 $[nedia] $X=46920 $Y=-4850 $dt=0
X5 2 3 4 1 LDDN w=5e-05 l=1.25e-06 adio=6.71697e-10 pdio=3.30958e-05 extlay=1 $[nedia] $X=58820 $Y=-4850 $dt=0
X6 2 3 4 1 LDDN w=5e-05 l=1.25e-06 adio=6.71697e-10 pdio=3.30958e-05 extlay=1 $[nedia] $X=70720 $Y=-4850 $dt=0
X7 2 3 4 1 LDDN w=5e-05 l=1.25e-06 adio=6.71697e-10 pdio=3.30958e-05 extlay=1 $[nedia] $X=82620 $Y=-4850 $dt=0
X8 2 3 4 1 LDDN w=5e-05 l=1.25e-06 adio=6.71697e-10 pdio=3.30958e-05 extlay=1 $[nedia] $X=94520 $Y=-4850 $dt=0
X9 2 3 4 1 LDDN w=5e-05 l=1.25e-06 adio=6.71697e-10 pdio=3.30958e-05 extlay=1 $[nedia] $X=106420 $Y=-4850 $dt=0
X10 2 3 4 1 LDDN w=5e-05 l=1.25e-06 adio=6.71697e-10 pdio=3.30958e-05 extlay=1 $[nedia] $X=118320 $Y=-4850 $dt=0
X11 2 3 4 1 LDDN w=5e-05 l=1.25e-06 adio=6.71697e-10 pdio=3.30958e-05 extlay=1 $[nedia] $X=130220 $Y=-4850 $dt=0
.ends nedia_CDNS_723062655410

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X12                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X12 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7230626554116 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7230626554116 $T=500 1500 0 0 $X=0 $Y=1000
X2 1 VIATP_C_CDNS_7230626554116 $T=500 2500 0 0 $X=0 $Y=2000
X3 1 VIATP_C_CDNS_7230626554116 $T=500 3500 0 0 $X=0 $Y=3000
X4 1 VIATP_C_CDNS_7230626554116 $T=500 4500 0 0 $X=0 $Y=4000
X5 1 VIATP_C_CDNS_7230626554116 $T=500 5500 0 0 $X=0 $Y=5000
X6 1 VIATP_C_CDNS_7230626554116 $T=500 6500 0 0 $X=0 $Y=6000
X7 1 VIATP_C_CDNS_7230626554116 $T=500 7500 0 0 $X=0 $Y=7000
X8 1 VIATP_C_CDNS_7230626554116 $T=500 8500 0 0 $X=0 $Y=8000
X9 1 VIATP_C_CDNS_7230626554116 $T=500 9500 0 0 $X=0 $Y=9000
.ends MASCO__X12

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X14                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X14 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7230626554116 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7230626554116 $T=500 2500 0 0 $X=0 $Y=2000
X2 1 VIATP_C_CDNS_7230626554116 $T=500 4500 0 0 $X=0 $Y=4000
X3 1 VIATP_C_CDNS_7230626554116 $T=500 6500 0 0 $X=0 $Y=6000
X4 1 VIATP_C_CDNS_7230626554116 $T=500 8500 0 0 $X=0 $Y=8000
.ends MASCO__X14

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y18                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y18 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7230626554136 $T=500 620 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7230626554136 $T=1500 620 0 0 $X=1000 $Y=0
X2 1 VIATP_C_CDNS_7230626554136 $T=2500 620 0 0 $X=2000 $Y=0
X3 1 VIATP_C_CDNS_7230626554136 $T=3500 620 0 0 $X=3000 $Y=0
X4 1 VIATP_C_CDNS_7230626554136 $T=4500 620 0 0 $X=4000 $Y=0
X5 1 VIATP_C_CDNS_7230626554136 $T=5500 620 0 0 $X=5000 $Y=0
X6 1 VIATP_C_CDNS_7230626554136 $T=6500 620 0 0 $X=6000 $Y=0
X7 1 VIATP_C_CDNS_7230626554136 $T=7500 620 0 0 $X=7000 $Y=0
X8 1 VIATP_C_CDNS_7230626554136 $T=8500 620 0 0 $X=8000 $Y=0
X9 1 VIATP_C_CDNS_7230626554136 $T=9500 620 0 0 $X=9000 $Y=0
X10 1 VIATP_C_CDNS_7230626554136 $T=10500 620 0 0 $X=10000 $Y=0
X11 1 VIATP_C_CDNS_7230626554136 $T=11500 620 0 0 $X=11000 $Y=0
.ends MASCO__Y18

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y25                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y25 1
** N=1 EP=1 FDC=0
X0 1 MASCO__X14 $T=0 0 0 0 $X=0 $Y=0
X1 1 MASCO__X14 $T=2000 0 0 0 $X=2000 $Y=0
X2 1 MASCO__X14 $T=4000 0 0 0 $X=4000 $Y=0
X3 1 MASCO__X14 $T=6000 0 0 0 $X=6000 $Y=0
X4 1 MASCO__X14 $T=8000 0 0 0 $X=8000 $Y=0
X5 1 MASCO__X14 $T=10000 0 0 0 $X=10000 $Y=0
X6 1 MASCO__X14 $T=12000 0 0 0 $X=12000 $Y=0
X7 1 MASCO__X14 $T=14000 0 0 0 $X=14000 $Y=0
.ends MASCO__Y25

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y26                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y26 1
** N=1 EP=1 FDC=0
X0 1 MASCO__X12 $T=0 0 0 0 $X=0 $Y=0
X1 1 MASCO__X12 $T=2000 0 0 0 $X=2000 $Y=0
X2 1 MASCO__X12 $T=4000 0 0 0 $X=4000 $Y=0
X3 1 MASCO__X12 $T=6000 0 0 0 $X=6000 $Y=0
X4 1 MASCO__X12 $T=8000 0 0 0 $X=8000 $Y=0
X5 1 MASCO__X12 $T=10000 0 0 0 $X=10000 $Y=0
X6 1 MASCO__X12 $T=12000 0 0 0 $X=12000 $Y=0
X7 1 MASCO__X12 $T=14000 0 0 0 $X=14000 $Y=0
.ends MASCO__Y26

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__H1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__H1 1 2 3 4
** N=4 EP=4 FDC=12
X0 4 VIATP_C_CDNS_7230626554116 $T=375420 65345 0 0 $X=374920 $Y=64845
X1 4 VIATP_C_CDNS_7230626554136 $T=263420 75465 0 0 $X=262920 $Y=74845
X2 3 VIATP_C_CDNS_7230626554136 $T=287035 117625 0 0 $X=286535 $Y=117005
X3 3 VIATP_C_CDNS_7230626554136 $T=288035 117625 0 0 $X=287535 $Y=117005
X4 3 VIATP_C_CDNS_7230626554136 $T=289035 117625 0 0 $X=288535 $Y=117005
X5 3 VIATP_C_CDNS_7230626554136 $T=290035 117625 0 0 $X=289535 $Y=117005
X6 3 VIATP_C_CDNS_7230626554136 $T=291035 117625 0 0 $X=290535 $Y=117005
X7 3 VIATP_C_CDNS_7230626554136 $T=292035 117625 0 0 $X=291535 $Y=117005
X8 3 VIATP_C_CDNS_7230626554136 $T=293035 117625 0 0 $X=292535 $Y=117005
X9 3 VIATP_C_CDNS_7230626554136 $T=294035 117625 0 0 $X=293535 $Y=117005
X10 3 VIATP_C_CDNS_7230626554136 $T=295035 117625 0 0 $X=294535 $Y=117005
X11 3 VIATP_C_CDNS_7230626554136 $T=296035 117625 0 0 $X=295535 $Y=117005
X12 4 VIATP_C_CDNS_7230626554136 $T=372420 75465 0 0 $X=371920 $Y=74845
X13 4 VIATP_C_CDNS_7230626554136 $T=373420 75465 0 0 $X=372920 $Y=74845
X14 4 VIATP_C_CDNS_7230626554136 $T=374420 75465 0 0 $X=373920 $Y=74845
X15 3 VIATP_C_CDNS_7230626554136 $T=395035 117625 0 0 $X=394535 $Y=117005
X16 3 VIATP_C_CDNS_7230626554136 $T=396035 117625 0 0 $X=395535 $Y=117005
X17 3 VIATP_C_CDNS_7230626554136 $T=397035 117625 0 0 $X=396535 $Y=117005
X18 3 VIATP_C_CDNS_7230626554136 $T=398035 117625 0 0 $X=397535 $Y=117005
X19 3 VIATP_C_CDNS_7230626554136 $T=399035 117625 0 0 $X=398535 $Y=117005
X20 3 VIATP_C_CDNS_7230626554136 $T=400035 117625 0 0 $X=399535 $Y=117005
X21 3 VIATP_C_CDNS_7230626554136 $T=401035 117625 0 0 $X=400535 $Y=117005
X22 4 VIATP_C_CDNS_7230626554136 $T=401420 75465 0 0 $X=400920 $Y=74845
X23 3 VIATP_C_CDNS_7230626554136 $T=402035 117625 0 0 $X=401535 $Y=117005
X24 4 VIATP_C_CDNS_7230626554136 $T=402420 75465 0 0 $X=401920 $Y=74845
X25 3 VIATP_C_CDNS_7230626554136 $T=403035 117625 0 0 $X=402535 $Y=117005
X26 4 VIATP_C_CDNS_7230626554136 $T=403420 75465 0 0 $X=402920 $Y=74845
X27 3 VIATP_C_CDNS_7230626554136 $T=404035 117625 0 0 $X=403535 $Y=117005
X28 4 VIATP_C_CDNS_7230626554136 $T=404420 75465 0 0 $X=403920 $Y=74845
X29 3 VIATP_C_CDNS_7230626554136 $T=405035 117625 0 0 $X=404535 $Y=117005
X30 4 VIATP_C_CDNS_7230626554136 $T=405420 75465 0 0 $X=404920 $Y=74845
X31 3 VIATP_C_CDNS_7230626554136 $T=407035 117625 0 0 $X=406535 $Y=117005
X32 4 VIATP_C_CDNS_7230626554136 $T=407420 75465 0 0 $X=406920 $Y=74845
X33 3 VIATP_C_CDNS_7230626554136 $T=408035 117625 0 0 $X=407535 $Y=117005
X34 4 VIATP_C_CDNS_7230626554136 $T=408420 75465 0 0 $X=407920 $Y=74845
X35 3 VIATP_C_CDNS_7230626554136 $T=409035 117625 0 0 $X=408535 $Y=117005
X36 4 VIATP_C_CDNS_7230626554136 $T=409420 75465 0 0 $X=408920 $Y=74845
X37 3 VIATP_C_CDNS_7230626554136 $T=410035 117625 0 0 $X=409535 $Y=117005
X38 4 VIATP_C_CDNS_7230626554136 $T=410420 75465 0 0 $X=409920 $Y=74845
X39 3 VIATP_C_CDNS_7230626554136 $T=411035 117625 0 0 $X=410535 $Y=117005
X40 4 VIATP_C_CDNS_7230626554136 $T=411420 75465 0 0 $X=410920 $Y=74845
X41 3 VIATP_C_CDNS_7230626554136 $T=412035 117625 0 0 $X=411535 $Y=117005
X42 4 VIATP_C_CDNS_7230626554136 $T=412420 75465 0 0 $X=411920 $Y=74845
X43 3 VIATP_C_CDNS_7230626554136 $T=413035 117625 0 0 $X=412535 $Y=117005
X44 4 VIATP_C_CDNS_7230626554136 $T=413420 75465 0 0 $X=412920 $Y=74845
X45 3 VIATP_C_CDNS_7230626554136 $T=414035 117625 0 0 $X=413535 $Y=117005
X46 4 VIATP_C_CDNS_7230626554136 $T=414420 75465 0 0 $X=413920 $Y=74845
X47 4 VIATP_C_CDNS_7230626554137 $T=406480 75465 0 0 $X=406040 $Y=74845
X48 3 VIATP_C_CDNS_7230626554145 $T=405785 118745 0 0 $X=405515 $Y=118245
X49 3 VIATP_C_CDNS_7230626554145 $T=405785 119745 0 0 $X=405515 $Y=119245
X50 3 VIATP_C_CDNS_7230626554145 $T=405785 120745 0 0 $X=405515 $Y=120245
X51 3 VIATP_C_CDNS_7230626554145 $T=405785 121745 0 0 $X=405515 $Y=121245
X52 3 VIATP_C_CDNS_7230626554145 $T=405785 122745 0 0 $X=405515 $Y=122245
X53 3 VIATP_C_CDNS_7230626554145 $T=405785 123745 0 0 $X=405515 $Y=123245
X54 3 VIATP_C_CDNS_7230626554145 $T=405785 124745 0 0 $X=405515 $Y=124245
X55 3 VIATP_C_CDNS_7230626554145 $T=405785 125745 0 0 $X=405515 $Y=125245
X56 3 VIATP_C_CDNS_7230626554145 $T=405785 126745 0 0 $X=405515 $Y=126245
X57 3 VIATP_C_CDNS_7230626554145 $T=405785 127745 0 0 $X=405515 $Y=127245
X58 3 VIATP_C_CDNS_7230626554149 $T=261795 117625 0 0 $X=261065 $Y=117005
X59 3 VIATP_C_CDNS_7230626554150 $T=297685 118745 0 0 $X=297415 $Y=118245
X60 3 VIATP_C_CDNS_7230626554150 $T=297685 119745 0 0 $X=297415 $Y=119245
X61 3 VIATP_C_CDNS_7230626554150 $T=297685 120745 0 0 $X=297415 $Y=120245
X62 3 VIATP_C_CDNS_7230626554150 $T=297685 121745 0 0 $X=297415 $Y=121245
X63 3 VIATP_C_CDNS_7230626554150 $T=297685 122745 0 0 $X=297415 $Y=122245
X64 3 VIATP_C_CDNS_7230626554150 $T=297685 123745 0 0 $X=297415 $Y=123245
X65 3 VIATP_C_CDNS_7230626554150 $T=297685 124745 0 0 $X=297415 $Y=124245
X66 3 VIATP_C_CDNS_7230626554150 $T=297685 125745 0 0 $X=297415 $Y=125245
X67 3 VIATP_C_CDNS_7230626554150 $T=297685 126745 0 0 $X=297415 $Y=126245
X68 3 VIATP_C_CDNS_7230626554150 $T=297685 127745 0 0 $X=297415 $Y=127245
X69 3 VIATP_C_CDNS_7230626554151 $T=261795 118745 0 0 $X=261065 $Y=118245
X70 3 VIATP_C_CDNS_7230626554151 $T=261795 119745 0 0 $X=261065 $Y=119245
X71 3 VIATP_C_CDNS_7230626554151 $T=261795 120745 0 0 $X=261065 $Y=120245
X72 3 VIATP_C_CDNS_7230626554151 $T=261795 121745 0 0 $X=261065 $Y=121245
X73 3 VIATP_C_CDNS_7230626554151 $T=261795 122745 0 0 $X=261065 $Y=122245
X74 3 VIATP_C_CDNS_7230626554151 $T=261795 123745 0 0 $X=261065 $Y=123245
X75 3 VIATP_C_CDNS_7230626554151 $T=261795 124745 0 0 $X=261065 $Y=124245
X76 3 VIATP_C_CDNS_7230626554151 $T=261795 125745 0 0 $X=261065 $Y=125245
X77 3 VIATP_C_CDNS_7230626554151 $T=261795 126745 0 0 $X=261065 $Y=126245
X78 3 VIATP_C_CDNS_7230626554151 $T=261795 127745 0 0 $X=261065 $Y=127245
X79 4 VIATP_C_CDNS_7230626554153 $T=261990 75465 0 0 $X=261060 $Y=74845
X80 4 VIATP_C_CDNS_7230626554154 $T=261990 65345 0 0 $X=261060 $Y=64845
X81 4 VIATP_C_CDNS_7230626554154 $T=261990 66345 0 0 $X=261060 $Y=65845
X82 4 VIATP_C_CDNS_7230626554154 $T=261990 67345 0 0 $X=261060 $Y=66845
X83 4 VIATP_C_CDNS_7230626554154 $T=261990 68345 0 0 $X=261060 $Y=67845
X84 4 VIATP_C_CDNS_7230626554154 $T=261990 69345 0 0 $X=261060 $Y=68845
X85 4 VIATP_C_CDNS_7230626554154 $T=261990 70345 0 0 $X=261060 $Y=69845
X86 4 VIATP_C_CDNS_7230626554154 $T=261990 71345 0 0 $X=261060 $Y=70845
X87 4 VIATP_C_CDNS_7230626554154 $T=261990 72345 0 0 $X=261060 $Y=71845
X88 4 VIATP_C_CDNS_7230626554154 $T=261990 73345 0 0 $X=261060 $Y=72845
X89 4 VIATP_C_CDNS_7230626554154 $T=261990 74345 0 0 $X=261060 $Y=73845
X90 4 VIATP_C_CDNS_7230626554157 $T=406480 65345 0 0 $X=406040 $Y=64845
X91 4 VIATP_C_CDNS_7230626554157 $T=406480 66345 0 0 $X=406040 $Y=65845
X92 4 VIATP_C_CDNS_7230626554157 $T=406480 67345 0 0 $X=406040 $Y=66845
X93 4 VIATP_C_CDNS_7230626554157 $T=406480 68345 0 0 $X=406040 $Y=67845
X94 4 VIATP_C_CDNS_7230626554157 $T=406480 69345 0 0 $X=406040 $Y=68845
X95 4 VIATP_C_CDNS_7230626554157 $T=406480 70345 0 0 $X=406040 $Y=69845
X96 4 VIATP_C_CDNS_7230626554157 $T=406480 71345 0 0 $X=406040 $Y=70845
X97 4 VIATP_C_CDNS_7230626554157 $T=406480 72345 0 0 $X=406040 $Y=71845
X98 4 VIATP_C_CDNS_7230626554157 $T=406480 73345 0 0 $X=406040 $Y=72845
X99 4 VIATP_C_CDNS_7230626554157 $T=406480 74345 0 0 $X=406040 $Y=73845
X100 4 VIATP_C_CDNS_7230626554158 $T=375550 67345 0 0 $X=375185 $Y=66845
X101 4 VIATP_C_CDNS_7230626554158 $T=375550 69345 0 0 $X=375185 $Y=68845
X102 4 VIATP_C_CDNS_7230626554158 $T=375550 71345 0 0 $X=375185 $Y=70845
X103 4 VIATP_C_CDNS_7230626554158 $T=375550 73345 0 0 $X=375185 $Y=72845
X104 1 3 2 4 nedia_CDNS_723062655410 $T=267970 84045 0 0 $X=251750 $Y=64655
X105 3 MASCO__X12 $T=263535 118245 0 0 $X=263535 $Y=118245
X106 3 MASCO__X12 $T=265535 118245 0 0 $X=265535 $Y=118245
X107 3 MASCO__X12 $T=267535 118245 0 0 $X=267535 $Y=118245
X108 3 MASCO__X12 $T=269535 118245 0 0 $X=269535 $Y=118245
X109 3 MASCO__X12 $T=271535 118245 0 0 $X=271535 $Y=118245
X110 3 MASCO__X12 $T=273535 118245 0 0 $X=273535 $Y=118245
X111 3 MASCO__X12 $T=275535 118245 0 0 $X=275535 $Y=118245
X112 3 MASCO__X12 $T=277535 118245 0 0 $X=277535 $Y=118245
X113 3 MASCO__X12 $T=279535 118245 0 0 $X=279535 $Y=118245
X114 3 MASCO__X12 $T=299535 118245 0 0 $X=299535 $Y=118245
X115 3 MASCO__X12 $T=301535 118245 0 0 $X=301535 $Y=118245
X116 3 MASCO__X12 $T=303535 118245 0 0 $X=303535 $Y=118245
X117 3 MASCO__X12 $T=305535 118245 0 0 $X=305535 $Y=118245
X118 3 MASCO__X12 $T=307535 118245 0 0 $X=307535 $Y=118245
X119 3 MASCO__X12 $T=309535 118245 0 0 $X=309535 $Y=118245
X120 3 MASCO__X12 $T=311535 118245 0 0 $X=311535 $Y=118245
X121 3 MASCO__X12 $T=313535 118245 0 0 $X=313535 $Y=118245
X122 3 MASCO__X12 $T=315535 118245 0 0 $X=315535 $Y=118245
X123 3 MASCO__X12 $T=317535 118245 0 0 $X=317535 $Y=118245
X124 3 MASCO__X12 $T=319535 118245 0 0 $X=319535 $Y=118245
X125 3 MASCO__X12 $T=321535 118245 0 0 $X=321535 $Y=118245
X126 3 MASCO__X12 $T=323535 118245 0 0 $X=323535 $Y=118245
X127 3 MASCO__X12 $T=325535 118245 0 0 $X=325535 $Y=118245
X128 3 MASCO__X12 $T=327535 118245 0 0 $X=327535 $Y=118245
X129 3 MASCO__X12 $T=329535 118245 0 0 $X=329535 $Y=118245
X130 3 MASCO__X12 $T=331535 118245 0 0 $X=331535 $Y=118245
X131 3 MASCO__X12 $T=333535 118245 0 0 $X=333535 $Y=118245
X132 3 MASCO__X12 $T=335535 118245 0 0 $X=335535 $Y=118245
X133 3 MASCO__X12 $T=337535 118245 0 0 $X=337535 $Y=118245
X134 3 MASCO__X12 $T=339535 118245 0 0 $X=339535 $Y=118245
X135 3 MASCO__X12 $T=341535 118245 0 0 $X=341535 $Y=118245
X136 3 MASCO__X12 $T=343535 118245 0 0 $X=343535 $Y=118245
X137 3 MASCO__X12 $T=345535 118245 0 0 $X=345535 $Y=118245
X138 3 MASCO__X12 $T=347535 118245 0 0 $X=347535 $Y=118245
X139 3 MASCO__X12 $T=349535 118245 0 0 $X=349535 $Y=118245
X140 3 MASCO__X12 $T=351535 118245 0 0 $X=351535 $Y=118245
X141 3 MASCO__X12 $T=353535 118245 0 0 $X=353535 $Y=118245
X142 3 MASCO__X12 $T=355535 118245 0 0 $X=355535 $Y=118245
X143 3 MASCO__X12 $T=357535 118245 0 0 $X=357535 $Y=118245
X144 3 MASCO__X12 $T=359535 118245 0 0 $X=359535 $Y=118245
X145 3 MASCO__X12 $T=361535 118245 0 0 $X=361535 $Y=118245
X146 3 MASCO__X12 $T=363535 118245 0 0 $X=363535 $Y=118245
X147 3 MASCO__X12 $T=365535 118245 0 0 $X=365535 $Y=118245
X148 3 MASCO__X12 $T=367535 118245 0 0 $X=367535 $Y=118245
X149 3 MASCO__X12 $T=369535 118245 0 0 $X=369535 $Y=118245
X150 3 MASCO__X12 $T=371535 118245 0 0 $X=371535 $Y=118245
X151 3 MASCO__X12 $T=373535 118245 0 0 $X=373535 $Y=118245
X152 3 MASCO__X12 $T=375535 118245 0 0 $X=375535 $Y=118245
X153 3 MASCO__X12 $T=377535 118245 0 0 $X=377535 $Y=118245
X154 4 MASCO__X12 $T=377920 64845 0 0 $X=377920 $Y=64845
X155 3 MASCO__X12 $T=379535 118245 0 0 $X=379535 $Y=118245
X156 4 MASCO__X12 $T=379920 64845 0 0 $X=379920 $Y=64845
X157 3 MASCO__X12 $T=381535 118245 0 0 $X=381535 $Y=118245
X158 4 MASCO__X12 $T=381920 64845 0 0 $X=381920 $Y=64845
X159 3 MASCO__X12 $T=383535 118245 0 0 $X=383535 $Y=118245
X160 4 MASCO__X12 $T=383920 64845 0 0 $X=383920 $Y=64845
X161 3 MASCO__X12 $T=385535 118245 0 0 $X=385535 $Y=118245
X162 4 MASCO__X12 $T=385920 64845 0 0 $X=385920 $Y=64845
X163 3 MASCO__X12 $T=387535 118245 0 0 $X=387535 $Y=118245
X164 4 MASCO__X12 $T=387920 64845 0 0 $X=387920 $Y=64845
X165 3 MASCO__X12 $T=389535 118245 0 0 $X=389535 $Y=118245
X166 4 MASCO__X12 $T=389920 64845 0 0 $X=389920 $Y=64845
X167 3 MASCO__X12 $T=391535 118245 0 0 $X=391535 $Y=118245
X168 4 MASCO__X12 $T=391920 64845 0 0 $X=391920 $Y=64845
X169 3 MASCO__X12 $T=393535 118245 0 0 $X=393535 $Y=118245
X170 4 MASCO__X12 $T=393920 64845 0 0 $X=393920 $Y=64845
X171 3 MASCO__X12 $T=395535 118245 0 0 $X=395535 $Y=118245
X172 4 MASCO__X12 $T=395920 64845 0 0 $X=395920 $Y=64845
X173 3 MASCO__X12 $T=397535 118245 0 0 $X=397535 $Y=118245
X174 4 MASCO__X12 $T=397920 64845 0 0 $X=397920 $Y=64845
X175 3 MASCO__X12 $T=399535 118245 0 0 $X=399535 $Y=118245
X176 4 MASCO__X12 $T=399920 64845 0 0 $X=399920 $Y=64845
X177 3 MASCO__X12 $T=401535 118245 0 0 $X=401535 $Y=118245
X178 4 MASCO__X12 $T=401920 64845 0 0 $X=401920 $Y=64845
X179 3 MASCO__X12 $T=403535 118245 0 0 $X=403535 $Y=118245
X180 4 MASCO__X12 $T=403920 64845 0 0 $X=403920 $Y=64845
X181 3 MASCO__X12 $T=407535 118245 0 0 $X=407535 $Y=118245
X182 4 MASCO__X12 $T=407920 64845 0 0 $X=407920 $Y=64845
X183 3 MASCO__X12 $T=409535 118245 0 0 $X=409535 $Y=118245
X184 4 MASCO__X12 $T=409920 64845 0 0 $X=409920 $Y=64845
X185 3 MASCO__X12 $T=411535 118245 0 0 $X=411535 $Y=118245
X186 4 MASCO__X12 $T=411920 64845 0 0 $X=411920 $Y=64845
X187 3 MASCO__X12 $T=413535 118245 0 0 $X=413535 $Y=118245
X188 4 MASCO__X12 $T=413920 64845 0 0 $X=413920 $Y=64845
X189 3 MASCO__X14 $T=262535 119245 0 0 $X=262535 $Y=119245
X190 3 MASCO__X14 $T=264535 119245 0 0 $X=264535 $Y=119245
X191 3 MASCO__X14 $T=266535 119245 0 0 $X=266535 $Y=119245
X192 3 MASCO__X14 $T=268535 119245 0 0 $X=268535 $Y=119245
X193 3 MASCO__X14 $T=270535 119245 0 0 $X=270535 $Y=119245
X194 3 MASCO__X14 $T=272535 119245 0 0 $X=272535 $Y=119245
X195 3 MASCO__X14 $T=274535 119245 0 0 $X=274535 $Y=119245
X196 3 MASCO__X14 $T=276535 119245 0 0 $X=276535 $Y=119245
X197 3 MASCO__X14 $T=278535 119245 0 0 $X=278535 $Y=119245
X198 3 MASCO__X14 $T=298535 119245 0 0 $X=298535 $Y=119245
X199 3 MASCO__X14 $T=300535 119245 0 0 $X=300535 $Y=119245
X200 3 MASCO__X14 $T=302535 119245 0 0 $X=302535 $Y=119245
X201 3 MASCO__X14 $T=304535 119245 0 0 $X=304535 $Y=119245
X202 3 MASCO__X14 $T=306535 119245 0 0 $X=306535 $Y=119245
X203 3 MASCO__X14 $T=308535 119245 0 0 $X=308535 $Y=119245
X204 3 MASCO__X14 $T=310535 119245 0 0 $X=310535 $Y=119245
X205 3 MASCO__X14 $T=312535 119245 0 0 $X=312535 $Y=119245
X206 3 MASCO__X14 $T=314535 119245 0 0 $X=314535 $Y=119245
X207 3 MASCO__X14 $T=316535 119245 0 0 $X=316535 $Y=119245
X208 3 MASCO__X14 $T=318535 119245 0 0 $X=318535 $Y=119245
X209 3 MASCO__X14 $T=320535 119245 0 0 $X=320535 $Y=119245
X210 3 MASCO__X14 $T=322535 119245 0 0 $X=322535 $Y=119245
X211 3 MASCO__X14 $T=324535 119245 0 0 $X=324535 $Y=119245
X212 3 MASCO__X14 $T=326535 119245 0 0 $X=326535 $Y=119245
X213 3 MASCO__X14 $T=328535 119245 0 0 $X=328535 $Y=119245
X214 3 MASCO__X14 $T=330535 119245 0 0 $X=330535 $Y=119245
X215 3 MASCO__X14 $T=332535 119245 0 0 $X=332535 $Y=119245
X216 3 MASCO__X14 $T=334535 119245 0 0 $X=334535 $Y=119245
X217 3 MASCO__X14 $T=336535 119245 0 0 $X=336535 $Y=119245
X218 3 MASCO__X14 $T=338535 119245 0 0 $X=338535 $Y=119245
X219 3 MASCO__X14 $T=340535 119245 0 0 $X=340535 $Y=119245
X220 3 MASCO__X14 $T=342535 119245 0 0 $X=342535 $Y=119245
X221 3 MASCO__X14 $T=344535 119245 0 0 $X=344535 $Y=119245
X222 3 MASCO__X14 $T=346535 119245 0 0 $X=346535 $Y=119245
X223 3 MASCO__X14 $T=348535 119245 0 0 $X=348535 $Y=119245
X224 3 MASCO__X14 $T=350535 119245 0 0 $X=350535 $Y=119245
X225 3 MASCO__X14 $T=352535 119245 0 0 $X=352535 $Y=119245
X226 3 MASCO__X14 $T=354535 119245 0 0 $X=354535 $Y=119245
X227 3 MASCO__X14 $T=356535 119245 0 0 $X=356535 $Y=119245
X228 3 MASCO__X14 $T=358535 119245 0 0 $X=358535 $Y=119245
X229 3 MASCO__X14 $T=360535 119245 0 0 $X=360535 $Y=119245
X230 3 MASCO__X14 $T=362535 119245 0 0 $X=362535 $Y=119245
X231 3 MASCO__X14 $T=364535 119245 0 0 $X=364535 $Y=119245
X232 3 MASCO__X14 $T=366535 119245 0 0 $X=366535 $Y=119245
X233 3 MASCO__X14 $T=368535 119245 0 0 $X=368535 $Y=119245
X234 3 MASCO__X14 $T=370535 119245 0 0 $X=370535 $Y=119245
X235 3 MASCO__X14 $T=372535 119245 0 0 $X=372535 $Y=119245
X236 3 MASCO__X14 $T=374535 119245 0 0 $X=374535 $Y=119245
X237 3 MASCO__X14 $T=376535 119245 0 0 $X=376535 $Y=119245
X238 4 MASCO__X14 $T=376920 64845 0 0 $X=376920 $Y=64845
X239 3 MASCO__X14 $T=378535 119245 0 0 $X=378535 $Y=119245
X240 4 MASCO__X14 $T=378920 64845 0 0 $X=378920 $Y=64845
X241 3 MASCO__X14 $T=380535 119245 0 0 $X=380535 $Y=119245
X242 4 MASCO__X14 $T=380920 64845 0 0 $X=380920 $Y=64845
X243 3 MASCO__X14 $T=382535 119245 0 0 $X=382535 $Y=119245
X244 4 MASCO__X14 $T=382920 64845 0 0 $X=382920 $Y=64845
X245 3 MASCO__X14 $T=384535 119245 0 0 $X=384535 $Y=119245
X246 4 MASCO__X14 $T=384920 64845 0 0 $X=384920 $Y=64845
X247 3 MASCO__X14 $T=386535 119245 0 0 $X=386535 $Y=119245
X248 4 MASCO__X14 $T=386920 64845 0 0 $X=386920 $Y=64845
X249 3 MASCO__X14 $T=388535 119245 0 0 $X=388535 $Y=119245
X250 4 MASCO__X14 $T=388920 64845 0 0 $X=388920 $Y=64845
X251 3 MASCO__X14 $T=390535 119245 0 0 $X=390535 $Y=119245
X252 4 MASCO__X14 $T=390920 64845 0 0 $X=390920 $Y=64845
X253 3 MASCO__X14 $T=392535 119245 0 0 $X=392535 $Y=119245
X254 4 MASCO__X14 $T=392920 64845 0 0 $X=392920 $Y=64845
X255 3 MASCO__X14 $T=394535 119245 0 0 $X=394535 $Y=119245
X256 4 MASCO__X14 $T=394920 64845 0 0 $X=394920 $Y=64845
X257 3 MASCO__X14 $T=396535 119245 0 0 $X=396535 $Y=119245
X258 4 MASCO__X14 $T=396920 64845 0 0 $X=396920 $Y=64845
X259 3 MASCO__X14 $T=398535 119245 0 0 $X=398535 $Y=119245
X260 4 MASCO__X14 $T=398920 64845 0 0 $X=398920 $Y=64845
X261 3 MASCO__X14 $T=400535 119245 0 0 $X=400535 $Y=119245
X262 4 MASCO__X14 $T=400920 64845 0 0 $X=400920 $Y=64845
X263 3 MASCO__X14 $T=402535 119245 0 0 $X=402535 $Y=119245
X264 4 MASCO__X14 $T=402920 64845 0 0 $X=402920 $Y=64845
X265 4 MASCO__X14 $T=404920 64845 0 0 $X=404920 $Y=64845
X266 3 MASCO__X14 $T=406535 119245 0 0 $X=406535 $Y=119245
X267 4 MASCO__X14 $T=406920 64845 0 0 $X=406920 $Y=64845
X268 3 MASCO__X14 $T=408535 119245 0 0 $X=408535 $Y=119245
X269 4 MASCO__X14 $T=408920 64845 0 0 $X=408920 $Y=64845
X270 3 MASCO__X14 $T=410535 119245 0 0 $X=410535 $Y=119245
X271 4 MASCO__X14 $T=410920 64845 0 0 $X=410920 $Y=64845
X272 3 MASCO__X14 $T=412535 119245 0 0 $X=412535 $Y=119245
X273 4 MASCO__X14 $T=412920 64845 0 0 $X=412920 $Y=64845
X274 3 MASCO__Y18 $T=262535 117005 0 0 $X=262535 $Y=117005
X275 4 MASCO__Y18 $T=263920 74845 0 0 $X=263920 $Y=74845
X276 3 MASCO__Y18 $T=274535 117005 0 0 $X=274535 $Y=117005
X277 4 MASCO__Y18 $T=275920 74845 0 0 $X=275920 $Y=74845
X278 4 MASCO__Y18 $T=287920 74845 0 0 $X=287920 $Y=74845
X279 3 MASCO__Y18 $T=298535 117005 0 0 $X=298535 $Y=117005
X280 4 MASCO__Y18 $T=299920 74845 0 0 $X=299920 $Y=74845
X281 3 MASCO__Y18 $T=310535 117005 0 0 $X=310535 $Y=117005
X282 4 MASCO__Y18 $T=311920 74845 0 0 $X=311920 $Y=74845
X283 3 MASCO__Y18 $T=322535 117005 0 0 $X=322535 $Y=117005
X284 4 MASCO__Y18 $T=323920 74845 0 0 $X=323920 $Y=74845
X285 3 MASCO__Y18 $T=334535 117005 0 0 $X=334535 $Y=117005
X286 4 MASCO__Y18 $T=335920 74845 0 0 $X=335920 $Y=74845
X287 3 MASCO__Y18 $T=346535 117005 0 0 $X=346535 $Y=117005
X288 4 MASCO__Y18 $T=347920 74845 0 0 $X=347920 $Y=74845
X289 3 MASCO__Y18 $T=358535 117005 0 0 $X=358535 $Y=117005
X290 4 MASCO__Y18 $T=359920 74845 0 0 $X=359920 $Y=74845
X291 3 MASCO__Y18 $T=370535 117005 0 0 $X=370535 $Y=117005
X292 4 MASCO__Y18 $T=376920 74845 0 0 $X=376920 $Y=74845
X293 3 MASCO__Y18 $T=382535 117005 0 0 $X=382535 $Y=117005
X294 4 MASCO__Y18 $T=388920 74845 0 0 $X=388920 $Y=74845
X295 4 MASCO__Y25 $T=262920 64845 0 0 $X=262920 $Y=64845
X296 4 MASCO__Y25 $T=278920 64845 0 0 $X=278920 $Y=64845
X297 3 MASCO__Y25 $T=280535 119245 0 0 $X=280535 $Y=119245
X298 4 MASCO__Y25 $T=294920 64845 0 0 $X=294920 $Y=64845
X299 4 MASCO__Y25 $T=310920 64845 0 0 $X=310920 $Y=64845
X300 4 MASCO__Y25 $T=326920 64845 0 0 $X=326920 $Y=64845
X301 4 MASCO__Y25 $T=342920 64845 0 0 $X=342920 $Y=64845
X302 4 MASCO__Y25 $T=358920 64845 0 0 $X=358920 $Y=64845
X303 4 MASCO__Y26 $T=263920 64845 0 0 $X=263920 $Y=64845
X304 4 MASCO__Y26 $T=279920 64845 0 0 $X=279920 $Y=64845
X305 3 MASCO__Y26 $T=281535 118245 0 0 $X=281535 $Y=118245
X306 4 MASCO__Y26 $T=295920 64845 0 0 $X=295920 $Y=64845
X307 4 MASCO__Y26 $T=311920 64845 0 0 $X=311920 $Y=64845
X308 4 MASCO__Y26 $T=327920 64845 0 0 $X=327920 $Y=64845
X309 4 MASCO__Y26 $T=343920 64845 0 0 $X=343920 $Y=64845
X310 4 MASCO__Y26 $T=359920 64845 0 0 $X=359920 $Y=64845
.ends MASCO__H1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_723062655415                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_723062655415 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_723062655415

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nedia_CDNS_723062655413                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nedia_CDNS_723062655413 1 2 3 4
** N=4 EP=4 FDC=1
X0 2 4 3 1 LDDN w=2e-05 l=1.25e-06 adio=7.56916e-10 pdio=0.00010535 extlay=1 $[nedia] $X=-680 $Y=-4850 $dt=0
.ends nedia_CDNS_723062655413

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__H2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__H2 1 2 3 4
** N=4 EP=4 FDC=1
X0 2 VIA2_C_CDNS_723062655415 $T=60995 110945 0 0 $X=60765 $Y=109935
X1 2 VIA2_C_CDNS_723062655415 $T=60995 130365 0 0 $X=60765 $Y=129355
X2 1 3 4 2 nedia_CDNS_723062655413 $T=60995 115655 0 0 $X=44775 $Y=96265
.ends MASCO__H2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__H3                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__H3 1 2 3 4 5
** N=5 EP=5 FDC=1
X0 2 VIA2_C_CDNS_723062655415 $T=101020 110945 0 0 $X=100790 $Y=109935
X1 2 VIA2_C_CDNS_723062655415 $T=101020 130365 0 0 $X=100790 $Y=129355
X2 1 3 4 2 nedia_CDNS_723062655413 $T=101020 115655 0 0 $X=84800 $Y=96265
.ends MASCO__H3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_723062655410                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_723062655410 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_723062655410

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_723062655411                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_723062655411 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_723062655411

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_723062655417                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_723062655417 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_723062655417

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7230626554123                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7230626554123 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7230626554123

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7230626554134                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7230626554134 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7230626554134

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7230626554155                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7230626554155 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7230626554155

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_723062655414                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_723062655414 1 2 3 4
** N=4 EP=4 FDC=1
M0 3 2 1 4 ne3 L=3.5e-07 W=2.2e-07 AD=1.984e-13 AS=1.984e-13 PD=1.88e-06 PS=1.88e-06 $X=0 $Y=0 $dt=2
.ends ne3_CDNS_723062655414

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: dsba_CDNS_723062655417                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt dsba_CDNS_723062655417 1 2 3
** N=623 EP=3 FDC=21
D0 1 2 p_dwhn AREA=6.69221e-10 PJ=0.00022132 perimeter=0.00022132 $X=-3330 $Y=-3970 $dt=6
D1 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=1390 $Y=1050 $dt=8
D2 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=5350 $Y=1050 $dt=8
D3 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=9310 $Y=1050 $dt=8
D4 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=13270 $Y=1050 $dt=8
D5 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=17230 $Y=1050 $dt=8
D6 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=21190 $Y=1050 $dt=8
D7 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=25150 $Y=1050 $dt=8
D8 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=29110 $Y=1050 $dt=8
D9 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=33070 $Y=1050 $dt=8
D10 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=37030 $Y=1050 $dt=8
D11 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=40990 $Y=1050 $dt=8
D12 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=44950 $Y=1050 $dt=8
D13 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=48910 $Y=1050 $dt=8
D14 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=52870 $Y=1050 $dt=8
D15 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=56830 $Y=1050 $dt=8
D16 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=60790 $Y=1050 $dt=8
D17 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=64750 $Y=1050 $dt=8
D18 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=68710 $Y=1050 $dt=8
D19 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=72670 $Y=1050 $dt=8
D20 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=76630 $Y=1050 $dt=8
.ends dsba_CDNS_723062655417

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7230626554110                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7230626554110 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
M0 3 2 1 1 pe3 L=3e-07 W=4.4e-07 AD=2.112e-13 AS=2.112e-13 PD=1.84e-06 PS=1.84e-06 $X=0 $Y=0 $dt=3
.ends pe3_CDNS_7230626554110

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X6                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X6 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7230626554116 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7230626554116 $T=500 2500 0 0 $X=0 $Y=2000
X2 1 VIATP_C_CDNS_7230626554116 $T=500 4500 0 0 $X=0 $Y=4000
X3 1 VIATP_C_CDNS_7230626554116 $T=500 6500 0 0 $X=0 $Y=6000
X4 1 VIATP_C_CDNS_7230626554116 $T=500 8500 0 0 $X=0 $Y=8000
X5 1 VIATP_C_CDNS_7230626554116 $T=500 10500 0 0 $X=0 $Y=10000
.ends MASCO__X6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X7                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X7 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7230626554116 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7230626554116 $T=500 2500 0 0 $X=0 $Y=2000
X2 1 VIATP_C_CDNS_7230626554116 $T=500 4500 0 0 $X=0 $Y=4000
X3 1 VIATP_C_CDNS_7230626554116 $T=500 6500 0 0 $X=0 $Y=6000
X4 1 VIATP_C_CDNS_7230626554116 $T=500 8500 0 0 $X=0 $Y=8000
X5 1 VIATP_C_CDNS_7230626554116 $T=500 10500 0 0 $X=0 $Y=10000
X6 1 VIATP_C_CDNS_7230626554116 $T=500 12500 0 0 $X=0 $Y=12000
.ends MASCO__X7

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X8                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X8 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7230626554116 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7230626554116 $T=500 1500 0 0 $X=0 $Y=1000
X2 1 VIATP_C_CDNS_7230626554116 $T=500 2500 0 0 $X=0 $Y=2000
X3 1 VIATP_C_CDNS_7230626554116 $T=500 3500 0 0 $X=0 $Y=3000
X4 1 VIATP_C_CDNS_7230626554116 $T=500 4500 0 0 $X=0 $Y=4000
X5 1 VIATP_C_CDNS_7230626554116 $T=500 5500 0 0 $X=0 $Y=5000
X6 1 VIATP_C_CDNS_7230626554116 $T=500 6500 0 0 $X=0 $Y=6000
X7 1 VIATP_C_CDNS_7230626554116 $T=500 7500 0 0 $X=0 $Y=7000
X8 1 VIATP_C_CDNS_7230626554116 $T=500 8500 0 0 $X=0 $Y=8000
.ends MASCO__X8

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X9                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X9 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7230626554116 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7230626554116 $T=500 1500 0 0 $X=0 $Y=1000
X2 1 VIATP_C_CDNS_7230626554116 $T=500 2500 0 0 $X=0 $Y=2000
X3 1 VIATP_C_CDNS_7230626554116 $T=500 3500 0 0 $X=0 $Y=3000
X4 1 VIATP_C_CDNS_7230626554116 $T=500 4500 0 0 $X=0 $Y=4000
X5 1 VIATP_C_CDNS_7230626554116 $T=500 5500 0 0 $X=0 $Y=5000
X6 1 VIATP_C_CDNS_7230626554116 $T=500 6500 0 0 $X=0 $Y=6000
X7 1 VIATP_C_CDNS_7230626554116 $T=500 7500 0 0 $X=0 $Y=7000
.ends MASCO__X9

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y22                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y22 1
** N=1 EP=1 FDC=0
X0 1 MASCO__X8 $T=0 0 0 0 $X=0 $Y=0
X1 1 MASCO__X8 $T=2000 0 0 0 $X=2000 $Y=0
X2 1 MASCO__X8 $T=4000 0 0 0 $X=4000 $Y=0
X3 1 MASCO__X8 $T=6000 0 0 0 $X=6000 $Y=0
X4 1 MASCO__X8 $T=8000 0 0 0 $X=8000 $Y=0
X5 1 MASCO__X8 $T=10000 0 0 0 $X=10000 $Y=0
X6 1 MASCO__X8 $T=12000 0 0 0 $X=12000 $Y=0
X7 1 MASCO__X8 $T=14000 0 0 0 $X=14000 $Y=0
.ends MASCO__Y22

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y23                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y23 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7230626554134 $T=500 750 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7230626554134 $T=1500 750 0 0 $X=1000 $Y=0
X2 1 VIATP_C_CDNS_7230626554134 $T=2500 750 0 0 $X=2000 $Y=0
X3 1 VIATP_C_CDNS_7230626554134 $T=3500 750 0 0 $X=3000 $Y=0
X4 1 VIATP_C_CDNS_7230626554134 $T=4500 750 0 0 $X=4000 $Y=0
X5 1 VIATP_C_CDNS_7230626554134 $T=5500 750 0 0 $X=5000 $Y=0
X6 1 VIATP_C_CDNS_7230626554134 $T=6500 750 0 0 $X=6000 $Y=0
X7 1 VIATP_C_CDNS_7230626554134 $T=7500 750 0 0 $X=7000 $Y=0
X8 1 VIATP_C_CDNS_7230626554134 $T=8500 750 0 0 $X=8000 $Y=0
X9 1 VIATP_C_CDNS_7230626554134 $T=9500 750 0 0 $X=9000 $Y=0
X10 1 VIATP_C_CDNS_7230626554134 $T=10500 750 0 0 $X=10000 $Y=0
X11 1 VIATP_C_CDNS_7230626554134 $T=11500 750 0 0 $X=11000 $Y=0
.ends MASCO__Y23

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X10                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X10 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7230626554116 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7230626554116 $T=500 2500 0 0 $X=0 $Y=2000
X2 1 VIATP_C_CDNS_7230626554116 $T=500 4500 0 0 $X=0 $Y=4000
X3 1 VIATP_C_CDNS_7230626554116 $T=500 6500 0 0 $X=0 $Y=6000
X4 1 VIATP_C_CDNS_7230626554116 $T=500 8500 0 0 $X=0 $Y=8000
X5 1 VIATP_C_CDNS_7230626554116 $T=500 10500 0 0 $X=0 $Y=10000
X6 1 VIATP_C_CDNS_7230626554116 $T=500 12500 0 0 $X=0 $Y=12000
X7 1 VIATP_C_CDNS_7230626554116 $T=500 14500 0 0 $X=0 $Y=14000
.ends MASCO__X10

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y24                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y24 1
** N=1 EP=1 FDC=0
X0 1 MASCO__X10 $T=0 0 0 0 $X=0 $Y=0
X1 1 MASCO__X10 $T=2000 0 0 0 $X=2000 $Y=0
X2 1 MASCO__X10 $T=4000 0 0 0 $X=4000 $Y=0
X3 1 MASCO__X10 $T=6000 0 0 0 $X=6000 $Y=0
.ends MASCO__Y24

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__P4                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__P4 1 2 3 4 5 6 7 8 9 10
+ 11 12
** N=13 EP=12 FDC=399
X0 8 VIA1_C_CDNS_723062655410 $T=50810 88930 0 0 $X=50320 $Y=88700
X1 13 VIA1_C_CDNS_723062655410 $T=54130 88930 0 0 $X=53640 $Y=88700
X2 11 VIA1_C_CDNS_723062655410 $T=57450 88930 0 0 $X=56960 $Y=88700
X3 7 VIA1_C_CDNS_723062655411 $T=49730 85790 0 0 $X=49500 $Y=85300
X4 7 VIA1_C_CDNS_723062655411 $T=49730 87980 0 0 $X=49500 $Y=87490
X5 8 VIA1_C_CDNS_723062655411 $T=50640 85220 0 0 $X=50410 $Y=84730
X6 10 VIA1_C_CDNS_723062655411 $T=53050 85780 0 0 $X=52820 $Y=85290
X7 10 VIA1_C_CDNS_723062655411 $T=53050 87980 0 0 $X=52820 $Y=87490
X8 13 VIA1_C_CDNS_723062655411 $T=53985 85210 0 0 $X=53755 $Y=84720
X9 13 VIA1_C_CDNS_723062655411 $T=56370 85780 0 0 $X=56140 $Y=85290
X10 13 VIA1_C_CDNS_723062655411 $T=56370 87980 0 0 $X=56140 $Y=87490
X11 11 VIA1_C_CDNS_723062655411 $T=57305 85210 0 0 $X=57075 $Y=84720
X12 11 VIA2_C_CDNS_723062655415 $T=57470 89830 0 0 $X=57240 $Y=88820
X13 4 VIA1_C_CDNS_723062655417 $T=150435 94590 0 0 $X=150205 $Y=86300
X14 4 VIA1_C_CDNS_723062655417 $T=154395 94590 0 0 $X=154165 $Y=86300
X15 4 VIA1_C_CDNS_723062655417 $T=158355 94590 0 0 $X=158125 $Y=86300
X16 4 VIA1_C_CDNS_723062655417 $T=162315 94590 0 0 $X=162085 $Y=86300
X17 4 VIA1_C_CDNS_723062655417 $T=166280 94590 0 0 $X=166050 $Y=86300
X18 4 VIA1_C_CDNS_723062655417 $T=170240 94590 0 0 $X=170010 $Y=86300
X19 4 VIA1_C_CDNS_723062655417 $T=174200 94590 0 0 $X=173970 $Y=86300
X20 4 VIA1_C_CDNS_723062655417 $T=178160 94590 0 0 $X=177930 $Y=86300
X21 4 VIA1_C_CDNS_723062655417 $T=182115 94590 0 0 $X=181885 $Y=86300
X22 4 VIA1_C_CDNS_723062655417 $T=186075 94590 0 0 $X=185845 $Y=86300
X23 4 VIA1_C_CDNS_723062655417 $T=190035 94590 0 0 $X=189805 $Y=86300
X24 4 VIA1_C_CDNS_723062655417 $T=193995 94590 0 0 $X=193765 $Y=86300
X25 4 VIA1_C_CDNS_723062655417 $T=197960 94590 0 0 $X=197730 $Y=86300
X26 4 VIA1_C_CDNS_723062655417 $T=201920 94590 0 0 $X=201690 $Y=86300
X27 4 VIA1_C_CDNS_723062655417 $T=205880 94590 0 0 $X=205650 $Y=86300
X28 4 VIA1_C_CDNS_723062655417 $T=209840 94590 0 0 $X=209610 $Y=86300
X29 4 VIA1_C_CDNS_723062655417 $T=213795 94590 0 0 $X=213565 $Y=86300
X30 4 VIA1_C_CDNS_723062655417 $T=217755 94590 0 0 $X=217525 $Y=86300
X31 4 VIA1_C_CDNS_723062655417 $T=221715 94590 0 0 $X=221485 $Y=86300
X32 4 VIA1_C_CDNS_723062655417 $T=225675 94590 0 0 $X=225445 $Y=86300
X33 7 VIA2_C_CDNS_7230626554123 $T=49730 87120 0 0 $X=49500 $Y=86630
X34 10 VIA2_C_CDNS_7230626554123 $T=53050 86195 0 0 $X=52820 $Y=85705
X35 12 VIATP_C_CDNS_7230626554134 $T=371420 47095 0 0 $X=370920 $Y=46345
X36 12 VIATP_C_CDNS_7230626554134 $T=372420 47095 0 0 $X=371920 $Y=46345
X37 12 VIATP_C_CDNS_7230626554134 $T=373420 47095 0 0 $X=372920 $Y=46345
X38 12 VIATP_C_CDNS_7230626554134 $T=374420 47095 0 0 $X=373920 $Y=46345
X39 12 VIATP_C_CDNS_7230626554134 $T=375420 47095 0 0 $X=374920 $Y=46345
X40 12 VIATP_C_CDNS_7230626554134 $T=401420 47095 0 0 $X=400920 $Y=46345
X41 12 VIATP_C_CDNS_7230626554134 $T=402420 47095 0 0 $X=401920 $Y=46345
X42 12 VIATP_C_CDNS_7230626554134 $T=403420 47095 0 0 $X=402920 $Y=46345
X43 12 VIATP_C_CDNS_7230626554134 $T=404420 47095 0 0 $X=403920 $Y=46345
X44 12 VIATP_C_CDNS_7230626554134 $T=405420 47095 0 0 $X=404920 $Y=46345
X45 12 VIATP_C_CDNS_7230626554134 $T=407420 47095 0 0 $X=406920 $Y=46345
X46 12 VIATP_C_CDNS_7230626554134 $T=408420 47095 0 0 $X=407920 $Y=46345
X47 12 VIATP_C_CDNS_7230626554134 $T=409420 47095 0 0 $X=408920 $Y=46345
X48 12 VIATP_C_CDNS_7230626554134 $T=410420 47095 0 0 $X=409920 $Y=46345
X49 12 VIATP_C_CDNS_7230626554134 $T=411420 47095 0 0 $X=410920 $Y=46345
X50 12 VIATP_C_CDNS_7230626554134 $T=412420 47095 0 0 $X=411920 $Y=46345
X51 12 VIATP_C_CDNS_7230626554134 $T=413420 47095 0 0 $X=412920 $Y=46345
X52 12 VIATP_C_CDNS_7230626554134 $T=414420 47095 0 0 $X=413920 $Y=46345
X53 12 VIATP_C_CDNS_7230626554134 $T=415420 47095 0 0 $X=414920 $Y=46345
X54 12 VIATP_C_CDNS_7230626554134 $T=416420 47095 0 0 $X=415920 $Y=46345
X55 12 VIATP_C_CDNS_7230626554134 $T=417420 47095 0 0 $X=416920 $Y=46345
X56 12 VIATP_C_CDNS_7230626554134 $T=418420 47095 0 0 $X=417920 $Y=46345
X57 12 VIATP_C_CDNS_7230626554134 $T=419420 47095 0 0 $X=418920 $Y=46345
X58 12 VIATP_C_CDNS_7230626554134 $T=420420 47095 0 0 $X=419920 $Y=46345
X59 12 VIATP_C_CDNS_7230626554134 $T=421420 47095 0 0 $X=420920 $Y=46345
X60 12 VIATP_C_CDNS_7230626554134 $T=422420 47095 0 0 $X=421920 $Y=46345
X61 12 VIATP_C_CDNS_7230626554134 $T=423420 47095 0 0 $X=422920 $Y=46345
X62 12 VIATP_C_CDNS_7230626554134 $T=424420 47095 0 0 $X=423920 $Y=46345
X63 12 VIATP_C_CDNS_7230626554134 $T=425420 47095 0 0 $X=424920 $Y=46345
X64 12 VIATP_C_CDNS_7230626554134 $T=426420 47095 0 0 $X=425920 $Y=46345
X65 12 VIATP_C_CDNS_7230626554134 $T=427420 47095 0 0 $X=426920 $Y=46345
X66 12 VIATP_C_CDNS_7230626554134 $T=428420 47095 0 0 $X=427920 $Y=46345
X67 12 VIATP_C_CDNS_7230626554134 $T=429420 47095 0 0 $X=428920 $Y=46345
X68 12 VIATP_C_CDNS_7230626554134 $T=430420 47095 0 0 $X=429920 $Y=46345
X69 12 VIATP_C_CDNS_7230626554134 $T=431420 47095 0 0 $X=430920 $Y=46345
X70 12 VIATP_C_CDNS_7230626554136 $T=415420 75465 0 0 $X=414920 $Y=74845
X71 12 VIATP_C_CDNS_7230626554136 $T=416420 75465 0 0 $X=415920 $Y=74845
X72 12 VIATP_C_CDNS_7230626554136 $T=417420 75465 0 0 $X=416920 $Y=74845
X73 12 VIATP_C_CDNS_7230626554136 $T=418420 75465 0 0 $X=417920 $Y=74845
X74 12 VIATP_C_CDNS_7230626554136 $T=419420 75465 0 0 $X=418920 $Y=74845
X75 12 VIATP_C_CDNS_7230626554136 $T=420420 75465 0 0 $X=419920 $Y=74845
X76 12 VIATP_C_CDNS_7230626554136 $T=421420 75465 0 0 $X=420920 $Y=74845
X77 12 VIATP_C_CDNS_7230626554136 $T=422420 75465 0 0 $X=421920 $Y=74845
X78 12 VIATP_C_CDNS_7230626554136 $T=423420 75465 0 0 $X=422920 $Y=74845
X79 12 VIATP_C_CDNS_7230626554136 $T=424420 75465 0 0 $X=423920 $Y=74845
X80 12 VIATP_C_CDNS_7230626554136 $T=425420 75465 0 0 $X=424920 $Y=74845
X81 12 VIATP_C_CDNS_7230626554136 $T=426420 75465 0 0 $X=425920 $Y=74845
X82 12 VIATP_C_CDNS_7230626554136 $T=427420 75465 0 0 $X=426920 $Y=74845
X83 12 VIATP_C_CDNS_7230626554136 $T=428420 75465 0 0 $X=427920 $Y=74845
X84 12 VIATP_C_CDNS_7230626554136 $T=429420 75465 0 0 $X=428920 $Y=74845
X85 12 VIATP_C_CDNS_7230626554136 $T=430420 75465 0 0 $X=429920 $Y=74845
X86 12 VIATP_C_CDNS_7230626554136 $T=431420 75465 0 0 $X=430920 $Y=74845
X87 12 VIATP_C_CDNS_7230626554153 $T=432850 75465 0 0 $X=431920 $Y=74845
X88 12 VIATP_C_CDNS_7230626554154 $T=261990 48345 0 0 $X=261060 $Y=47845
X89 12 VIATP_C_CDNS_7230626554154 $T=261990 49345 0 0 $X=261060 $Y=48845
X90 12 VIATP_C_CDNS_7230626554154 $T=261990 50345 0 0 $X=261060 $Y=49845
X91 12 VIATP_C_CDNS_7230626554154 $T=261990 51345 0 0 $X=261060 $Y=50845
X92 12 VIATP_C_CDNS_7230626554154 $T=261990 52345 0 0 $X=261060 $Y=51845
X93 12 VIATP_C_CDNS_7230626554154 $T=261990 53345 0 0 $X=261060 $Y=52845
X94 12 VIATP_C_CDNS_7230626554154 $T=261990 54345 0 0 $X=261060 $Y=53845
X95 12 VIATP_C_CDNS_7230626554154 $T=261990 55345 0 0 $X=261060 $Y=54845
X96 12 VIATP_C_CDNS_7230626554154 $T=261990 56345 0 0 $X=261060 $Y=55845
X97 12 VIATP_C_CDNS_7230626554154 $T=261990 57345 0 0 $X=261060 $Y=56845
X98 12 VIATP_C_CDNS_7230626554154 $T=261990 58345 0 0 $X=261060 $Y=57845
X99 12 VIATP_C_CDNS_7230626554154 $T=261990 59345 0 0 $X=261060 $Y=58845
X100 12 VIATP_C_CDNS_7230626554154 $T=261990 60345 0 0 $X=261060 $Y=59845
X101 12 VIATP_C_CDNS_7230626554154 $T=261990 61345 0 0 $X=261060 $Y=60845
X102 12 VIATP_C_CDNS_7230626554154 $T=261990 62345 0 0 $X=261060 $Y=61845
X103 12 VIATP_C_CDNS_7230626554154 $T=261990 63345 0 0 $X=261060 $Y=62845
X104 12 VIATP_C_CDNS_7230626554154 $T=261990 64345 0 0 $X=261060 $Y=63845
X105 12 VIATP_C_CDNS_7230626554154 $T=432850 48345 0 0 $X=431920 $Y=47845
X106 12 VIATP_C_CDNS_7230626554154 $T=432850 49345 0 0 $X=431920 $Y=48845
X107 12 VIATP_C_CDNS_7230626554154 $T=432850 50345 0 0 $X=431920 $Y=49845
X108 12 VIATP_C_CDNS_7230626554154 $T=432850 51345 0 0 $X=431920 $Y=50845
X109 12 VIATP_C_CDNS_7230626554154 $T=432850 52345 0 0 $X=431920 $Y=51845
X110 12 VIATP_C_CDNS_7230626554154 $T=432850 53345 0 0 $X=431920 $Y=52845
X111 12 VIATP_C_CDNS_7230626554154 $T=432850 54345 0 0 $X=431920 $Y=53845
X112 12 VIATP_C_CDNS_7230626554154 $T=432850 55345 0 0 $X=431920 $Y=54845
X113 12 VIATP_C_CDNS_7230626554154 $T=432850 56345 0 0 $X=431920 $Y=55845
X114 12 VIATP_C_CDNS_7230626554154 $T=432850 57345 0 0 $X=431920 $Y=56845
X115 12 VIATP_C_CDNS_7230626554154 $T=432850 58345 0 0 $X=431920 $Y=57845
X116 12 VIATP_C_CDNS_7230626554154 $T=432850 59345 0 0 $X=431920 $Y=58845
X117 12 VIATP_C_CDNS_7230626554154 $T=432850 60345 0 0 $X=431920 $Y=59845
X118 12 VIATP_C_CDNS_7230626554154 $T=432850 61345 0 0 $X=431920 $Y=60845
X119 12 VIATP_C_CDNS_7230626554154 $T=432850 62345 0 0 $X=431920 $Y=61845
X120 12 VIATP_C_CDNS_7230626554154 $T=432850 63345 0 0 $X=431920 $Y=62845
X121 12 VIATP_C_CDNS_7230626554154 $T=432850 64345 0 0 $X=431920 $Y=63845
X122 12 VIATP_C_CDNS_7230626554154 $T=432850 65345 0 0 $X=431920 $Y=64845
X123 12 VIATP_C_CDNS_7230626554154 $T=432850 66345 0 0 $X=431920 $Y=65845
X124 12 VIATP_C_CDNS_7230626554154 $T=432850 67345 0 0 $X=431920 $Y=66845
X125 12 VIATP_C_CDNS_7230626554154 $T=432850 68345 0 0 $X=431920 $Y=67845
X126 12 VIATP_C_CDNS_7230626554154 $T=432850 69345 0 0 $X=431920 $Y=68845
X127 12 VIATP_C_CDNS_7230626554154 $T=432850 70345 0 0 $X=431920 $Y=69845
X128 12 VIATP_C_CDNS_7230626554154 $T=432850 71345 0 0 $X=431920 $Y=70845
X129 12 VIATP_C_CDNS_7230626554154 $T=432850 72345 0 0 $X=431920 $Y=71845
X130 12 VIATP_C_CDNS_7230626554154 $T=432850 73345 0 0 $X=431920 $Y=72845
X131 12 VIATP_C_CDNS_7230626554154 $T=432850 74345 0 0 $X=431920 $Y=73845
X132 12 VIATP_C_CDNS_7230626554155 $T=261990 47095 0 0 $X=261060 $Y=46345
X133 12 VIATP_C_CDNS_7230626554155 $T=432850 47095 0 0 $X=431920 $Y=46345
X134 12 VIATP_C_CDNS_7230626554157 $T=406480 48345 0 0 $X=406040 $Y=47845
X135 12 VIATP_C_CDNS_7230626554157 $T=406480 49345 0 0 $X=406040 $Y=48845
X136 12 VIATP_C_CDNS_7230626554157 $T=406480 50345 0 0 $X=406040 $Y=49845
X137 12 VIATP_C_CDNS_7230626554157 $T=406480 51345 0 0 $X=406040 $Y=50845
X138 12 VIATP_C_CDNS_7230626554157 $T=406480 52345 0 0 $X=406040 $Y=51845
X139 12 VIATP_C_CDNS_7230626554157 $T=406480 53345 0 0 $X=406040 $Y=52845
X140 12 VIATP_C_CDNS_7230626554157 $T=406480 54345 0 0 $X=406040 $Y=53845
X141 12 VIATP_C_CDNS_7230626554157 $T=406480 55345 0 0 $X=406040 $Y=54845
X142 12 VIATP_C_CDNS_7230626554157 $T=406480 56345 0 0 $X=406040 $Y=55845
X143 12 VIATP_C_CDNS_7230626554157 $T=406480 57345 0 0 $X=406040 $Y=56845
X144 12 VIATP_C_CDNS_7230626554157 $T=406480 58345 0 0 $X=406040 $Y=57845
X145 12 VIATP_C_CDNS_7230626554157 $T=406480 59345 0 0 $X=406040 $Y=58845
X146 12 VIATP_C_CDNS_7230626554157 $T=406480 60345 0 0 $X=406040 $Y=59845
X147 12 VIATP_C_CDNS_7230626554157 $T=406480 61345 0 0 $X=406040 $Y=60845
X148 12 VIATP_C_CDNS_7230626554157 $T=406480 62345 0 0 $X=406040 $Y=61845
X149 12 VIATP_C_CDNS_7230626554157 $T=406480 63345 0 0 $X=406040 $Y=62845
X150 12 VIATP_C_CDNS_7230626554157 $T=406480 64345 0 0 $X=406040 $Y=63845
X151 9 7 8 5 ne3_CDNS_723062655414 $T=49580 84790 0 0 $X=48740 $Y=84370
X152 9 10 13 5 ne3_CDNS_723062655414 $T=52925 84780 0 0 $X=52085 $Y=84360
X153 9 13 11 5 ne3_CDNS_723062655414 $T=56245 84780 0 0 $X=55405 $Y=84360
X154 5 3 4 dsba_CDNS_723062655417 $T=148575 85800 0 0 $X=140465 $Y=77050
X155 6 7 8 5 pe3_CDNS_7230626554110 $T=49580 89100 1 0 $X=48070 $Y=87630
X156 6 10 13 5 pe3_CDNS_7230626554110 $T=52900 89100 1 0 $X=51390 $Y=87630
X157 6 13 11 5 pe3_CDNS_7230626554110 $T=56220 89100 1 0 $X=54710 $Y=87630
X158 12 MASCO__X6 $T=414920 62845 0 0 $X=414920 $Y=62845
X159 12 MASCO__X6 $T=416920 62845 0 0 $X=416920 $Y=62845
X160 12 MASCO__X6 $T=418920 62845 0 0 $X=418920 $Y=62845
X161 12 MASCO__X6 $T=420920 62845 0 0 $X=420920 $Y=62845
X162 12 MASCO__X6 $T=422920 62845 0 0 $X=422920 $Y=62845
X163 12 MASCO__X6 $T=424920 62845 0 0 $X=424920 $Y=62845
X164 12 MASCO__X6 $T=426920 62845 0 0 $X=426920 $Y=62845
X165 12 MASCO__X6 $T=428920 62845 0 0 $X=428920 $Y=62845
X166 12 MASCO__X6 $T=430920 62845 0 0 $X=430920 $Y=62845
X167 12 MASCO__X7 $T=414920 48845 0 0 $X=414920 $Y=48845
X168 12 MASCO__X7 $T=416920 48845 0 0 $X=416920 $Y=48845
X169 12 MASCO__X7 $T=418920 48845 0 0 $X=418920 $Y=48845
X170 12 MASCO__X7 $T=420920 48845 0 0 $X=420920 $Y=48845
X171 12 MASCO__X7 $T=422920 48845 0 0 $X=422920 $Y=48845
X172 12 MASCO__X7 $T=424920 48845 0 0 $X=424920 $Y=48845
X173 12 MASCO__X7 $T=426920 48845 0 0 $X=426920 $Y=48845
X174 12 MASCO__X7 $T=428920 48845 0 0 $X=428920 $Y=48845
X175 12 MASCO__X7 $T=430920 48845 0 0 $X=430920 $Y=48845
X176 12 MASCO__X8 $T=377920 47845 0 0 $X=377920 $Y=47845
X177 12 MASCO__X8 $T=379920 47845 0 0 $X=379920 $Y=47845
X178 12 MASCO__X8 $T=381920 47845 0 0 $X=381920 $Y=47845
X179 12 MASCO__X8 $T=383920 47845 0 0 $X=383920 $Y=47845
X180 12 MASCO__X8 $T=385920 47845 0 0 $X=385920 $Y=47845
X181 12 MASCO__X8 $T=387920 47845 0 0 $X=387920 $Y=47845
X182 12 MASCO__X8 $T=389920 47845 0 0 $X=389920 $Y=47845
X183 12 MASCO__X8 $T=391920 47845 0 0 $X=391920 $Y=47845
X184 12 MASCO__X8 $T=393920 47845 0 0 $X=393920 $Y=47845
X185 12 MASCO__X8 $T=395920 47845 0 0 $X=395920 $Y=47845
X186 12 MASCO__X8 $T=397920 47845 0 0 $X=397920 $Y=47845
X187 12 MASCO__X8 $T=399920 47845 0 0 $X=399920 $Y=47845
X188 12 MASCO__X8 $T=401920 47845 0 0 $X=401920 $Y=47845
X189 12 MASCO__X8 $T=403920 47845 0 0 $X=403920 $Y=47845
X190 12 MASCO__X8 $T=407920 47845 0 0 $X=407920 $Y=47845
X191 12 MASCO__X8 $T=409920 47845 0 0 $X=409920 $Y=47845
X192 12 MASCO__X8 $T=411920 47845 0 0 $X=411920 $Y=47845
X193 12 MASCO__X8 $T=413920 47845 0 0 $X=413920 $Y=47845
X194 12 MASCO__X8 $T=415920 47845 0 0 $X=415920 $Y=47845
X195 12 MASCO__X8 $T=417920 47845 0 0 $X=417920 $Y=47845
X196 12 MASCO__X8 $T=419920 47845 0 0 $X=419920 $Y=47845
X197 12 MASCO__X8 $T=421920 47845 0 0 $X=421920 $Y=47845
X198 12 MASCO__X8 $T=423920 47845 0 0 $X=423920 $Y=47845
X199 12 MASCO__X8 $T=425920 47845 0 0 $X=425920 $Y=47845
X200 12 MASCO__X8 $T=427920 47845 0 0 $X=427920 $Y=47845
X201 12 MASCO__X8 $T=429920 47845 0 0 $X=429920 $Y=47845
X202 12 MASCO__X9 $T=263920 56845 0 0 $X=263920 $Y=56845
X203 12 MASCO__X9 $T=265920 56845 0 0 $X=265920 $Y=56845
X204 12 MASCO__X9 $T=267920 56845 0 0 $X=267920 $Y=56845
X205 12 MASCO__X9 $T=269920 56845 0 0 $X=269920 $Y=56845
X206 12 MASCO__X9 $T=271920 56845 0 0 $X=271920 $Y=56845
X207 12 MASCO__X9 $T=273920 56845 0 0 $X=273920 $Y=56845
X208 12 MASCO__X9 $T=275920 56845 0 0 $X=275920 $Y=56845
X209 12 MASCO__X9 $T=277920 56845 0 0 $X=277920 $Y=56845
X210 12 MASCO__X9 $T=279920 56845 0 0 $X=279920 $Y=56845
X211 12 MASCO__X9 $T=281920 56845 0 0 $X=281920 $Y=56845
X212 12 MASCO__X9 $T=283920 56845 0 0 $X=283920 $Y=56845
X213 12 MASCO__X9 $T=285920 56845 0 0 $X=285920 $Y=56845
X214 12 MASCO__X9 $T=287920 56845 0 0 $X=287920 $Y=56845
X215 12 MASCO__X9 $T=289920 56845 0 0 $X=289920 $Y=56845
X216 12 MASCO__X9 $T=291920 56845 0 0 $X=291920 $Y=56845
X217 12 MASCO__X9 $T=293920 56845 0 0 $X=293920 $Y=56845
X218 12 MASCO__X9 $T=295920 56845 0 0 $X=295920 $Y=56845
X219 12 MASCO__X9 $T=297920 56845 0 0 $X=297920 $Y=56845
X220 12 MASCO__X9 $T=299920 56845 0 0 $X=299920 $Y=56845
X221 12 MASCO__X9 $T=301920 56845 0 0 $X=301920 $Y=56845
X222 12 MASCO__X9 $T=303920 56845 0 0 $X=303920 $Y=56845
X223 12 MASCO__X9 $T=305920 56845 0 0 $X=305920 $Y=56845
X224 12 MASCO__X9 $T=307920 56845 0 0 $X=307920 $Y=56845
X225 12 MASCO__X9 $T=309920 56845 0 0 $X=309920 $Y=56845
X226 12 MASCO__X9 $T=311920 56845 0 0 $X=311920 $Y=56845
X227 12 MASCO__X9 $T=313920 56845 0 0 $X=313920 $Y=56845
X228 12 MASCO__X9 $T=315920 56845 0 0 $X=315920 $Y=56845
X229 12 MASCO__X9 $T=317920 56845 0 0 $X=317920 $Y=56845
X230 12 MASCO__X9 $T=319920 56845 0 0 $X=319920 $Y=56845
X231 12 MASCO__X9 $T=321920 56845 0 0 $X=321920 $Y=56845
X232 12 MASCO__X9 $T=323920 56845 0 0 $X=323920 $Y=56845
X233 12 MASCO__X9 $T=325920 56845 0 0 $X=325920 $Y=56845
X234 12 MASCO__X9 $T=327920 56845 0 0 $X=327920 $Y=56845
X235 12 MASCO__X9 $T=329920 56845 0 0 $X=329920 $Y=56845
X236 12 MASCO__X9 $T=331920 56845 0 0 $X=331920 $Y=56845
X237 12 MASCO__X9 $T=333920 56845 0 0 $X=333920 $Y=56845
X238 12 MASCO__X9 $T=335920 56845 0 0 $X=335920 $Y=56845
X239 12 MASCO__X9 $T=337920 56845 0 0 $X=337920 $Y=56845
X240 12 MASCO__X9 $T=339920 56845 0 0 $X=339920 $Y=56845
X241 12 MASCO__X9 $T=341920 56845 0 0 $X=341920 $Y=56845
X242 12 MASCO__X9 $T=343920 56845 0 0 $X=343920 $Y=56845
X243 12 MASCO__X9 $T=345920 56845 0 0 $X=345920 $Y=56845
X244 12 MASCO__X9 $T=347920 56845 0 0 $X=347920 $Y=56845
X245 12 MASCO__X9 $T=349920 56845 0 0 $X=349920 $Y=56845
X246 12 MASCO__X9 $T=351920 56845 0 0 $X=351920 $Y=56845
X247 12 MASCO__X9 $T=353920 56845 0 0 $X=353920 $Y=56845
X248 12 MASCO__X9 $T=355920 56845 0 0 $X=355920 $Y=56845
X249 12 MASCO__X9 $T=357920 56845 0 0 $X=357920 $Y=56845
X250 12 MASCO__X9 $T=359920 56845 0 0 $X=359920 $Y=56845
X251 12 MASCO__X9 $T=361920 56845 0 0 $X=361920 $Y=56845
X252 12 MASCO__X9 $T=363920 56845 0 0 $X=363920 $Y=56845
X253 12 MASCO__X9 $T=365920 56845 0 0 $X=365920 $Y=56845
X254 12 MASCO__X9 $T=367920 56845 0 0 $X=367920 $Y=56845
X255 12 MASCO__X9 $T=369920 56845 0 0 $X=369920 $Y=56845
X256 12 MASCO__X9 $T=371920 56845 0 0 $X=371920 $Y=56845
X257 12 MASCO__X9 $T=373920 56845 0 0 $X=373920 $Y=56845
X258 12 MASCO__X9 $T=377920 56845 0 0 $X=377920 $Y=56845
X259 12 MASCO__X9 $T=379920 56845 0 0 $X=379920 $Y=56845
X260 12 MASCO__X9 $T=381920 56845 0 0 $X=381920 $Y=56845
X261 12 MASCO__X9 $T=383920 56845 0 0 $X=383920 $Y=56845
X262 12 MASCO__X9 $T=385920 56845 0 0 $X=385920 $Y=56845
X263 12 MASCO__X9 $T=387920 56845 0 0 $X=387920 $Y=56845
X264 12 MASCO__X9 $T=389920 56845 0 0 $X=389920 $Y=56845
X265 12 MASCO__X9 $T=391920 56845 0 0 $X=391920 $Y=56845
X266 12 MASCO__X9 $T=393920 56845 0 0 $X=393920 $Y=56845
X267 12 MASCO__X9 $T=395920 56845 0 0 $X=395920 $Y=56845
X268 12 MASCO__X9 $T=397920 56845 0 0 $X=397920 $Y=56845
X269 12 MASCO__X9 $T=399920 56845 0 0 $X=399920 $Y=56845
X270 12 MASCO__X9 $T=401920 56845 0 0 $X=401920 $Y=56845
X271 12 MASCO__X9 $T=403920 56845 0 0 $X=403920 $Y=56845
X272 12 MASCO__X9 $T=407920 56845 0 0 $X=407920 $Y=56845
X273 12 MASCO__X9 $T=409920 56845 0 0 $X=409920 $Y=56845
X274 12 MASCO__X9 $T=411920 56845 0 0 $X=411920 $Y=56845
X275 12 MASCO__X9 $T=413920 56845 0 0 $X=413920 $Y=56845
X276 12 MASCO__Y22 $T=263920 47845 0 0 $X=263920 $Y=47845
X277 12 MASCO__Y22 $T=279920 47845 0 0 $X=279920 $Y=47845
X278 12 MASCO__Y22 $T=295920 47845 0 0 $X=295920 $Y=47845
X279 12 MASCO__Y22 $T=311920 47845 0 0 $X=311920 $Y=47845
X280 12 MASCO__Y22 $T=327920 47845 0 0 $X=327920 $Y=47845
X281 12 MASCO__Y22 $T=343920 47845 0 0 $X=343920 $Y=47845
X282 12 MASCO__Y22 $T=359920 47845 0 0 $X=359920 $Y=47845
X283 12 MASCO__Y22 $T=415920 56845 0 0 $X=415920 $Y=56845
X284 12 MASCO__Y22 $T=415920 65845 0 0 $X=415920 $Y=65845
X285 12 MASCO__Y23 $T=262920 46345 0 0 $X=262920 $Y=46345
X286 12 MASCO__Y23 $T=274920 46345 0 0 $X=274920 $Y=46345
X287 12 MASCO__Y23 $T=286920 46345 0 0 $X=286920 $Y=46345
X288 12 MASCO__Y23 $T=298920 46345 0 0 $X=298920 $Y=46345
X289 12 MASCO__Y23 $T=310920 46345 0 0 $X=310920 $Y=46345
X290 12 MASCO__Y23 $T=322920 46345 0 0 $X=322920 $Y=46345
X291 12 MASCO__Y23 $T=334920 46345 0 0 $X=334920 $Y=46345
X292 12 MASCO__Y23 $T=346920 46345 0 0 $X=346920 $Y=46345
X293 12 MASCO__Y23 $T=358920 46345 0 0 $X=358920 $Y=46345
X294 12 MASCO__Y23 $T=376920 46345 0 0 $X=376920 $Y=46345
X295 12 MASCO__Y23 $T=388920 46345 0 0 $X=388920 $Y=46345
X296 12 MASCO__Y24 $T=262920 48845 0 0 $X=262920 $Y=48845
X297 12 MASCO__Y24 $T=270920 48845 0 0 $X=270920 $Y=48845
X298 12 MASCO__Y24 $T=278920 48845 0 0 $X=278920 $Y=48845
X299 12 MASCO__Y24 $T=286920 48845 0 0 $X=286920 $Y=48845
X300 12 MASCO__Y24 $T=294920 48845 0 0 $X=294920 $Y=48845
X301 12 MASCO__Y24 $T=302920 48845 0 0 $X=302920 $Y=48845
X302 12 MASCO__Y24 $T=310920 48845 0 0 $X=310920 $Y=48845
X303 12 MASCO__Y24 $T=318920 48845 0 0 $X=318920 $Y=48845
X304 12 MASCO__Y24 $T=326920 48845 0 0 $X=326920 $Y=48845
X305 12 MASCO__Y24 $T=334920 48845 0 0 $X=334920 $Y=48845
X306 12 MASCO__Y24 $T=342920 48845 0 0 $X=342920 $Y=48845
X307 12 MASCO__Y24 $T=350920 48845 0 0 $X=350920 $Y=48845
X308 12 MASCO__Y24 $T=358920 48845 0 0 $X=358920 $Y=48845
X309 12 MASCO__Y24 $T=366920 48845 0 0 $X=366920 $Y=48845
X310 12 MASCO__Y24 $T=374920 48845 0 0 $X=374920 $Y=48845
X311 12 MASCO__Y24 $T=382920 48845 0 0 $X=382920 $Y=48845
X312 12 MASCO__Y24 $T=390920 48845 0 0 $X=390920 $Y=48845
X313 12 MASCO__Y24 $T=398920 48845 0 0 $X=398920 $Y=48845
X314 12 MASCO__Y24 $T=406920 48845 0 0 $X=406920 $Y=48845
D0 5 6 p_dnw AREA=3.39001e-11 PJ=3.421e-05 perimeter=3.421e-05 $X=46855 $Y=86465 $dt=4
D1 5 6 p_dnw3 AREA=2.49e-11 PJ=0 perimeter=0 $X=48070 $Y=87630 $dt=9
C2 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=-25270 $Y=-20340 $dt=11
C3 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=-25270 $Y=-8640 $dt=11
C4 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=-19230 $Y=-20340 $dt=11
C5 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=-19230 $Y=-8640 $dt=11
C6 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=-13190 $Y=-20340 $dt=11
C7 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=-13190 $Y=-8640 $dt=11
C8 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=-7150 $Y=-20340 $dt=11
C9 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=-7150 $Y=-8640 $dt=11
C10 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=-1110 $Y=-20340 $dt=11
C11 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=-1110 $Y=-8640 $dt=11
C12 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=4930 $Y=-20340 $dt=11
C13 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=4930 $Y=-8640 $dt=11
C14 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=10970 $Y=-20340 $dt=11
C15 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=10970 $Y=-8640 $dt=11
C16 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=17010 $Y=-20340 $dt=11
C17 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=17010 $Y=-8640 $dt=11
C18 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=23050 $Y=-20340 $dt=11
C19 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=23050 $Y=-8640 $dt=11
C20 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=29090 $Y=-20340 $dt=11
C21 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=29090 $Y=-8640 $dt=11
C22 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=35130 $Y=-20340 $dt=11
C23 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=35130 $Y=-8640 $dt=11
C24 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=40195 $Y=14580 $dt=11
C25 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=40195 $Y=20620 $dt=11
C26 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=40195 $Y=26660 $dt=11
C27 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=40195 $Y=32700 $dt=11
C28 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=40195 $Y=38740 $dt=11
C29 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=40195 $Y=44780 $dt=11
C30 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=40195 $Y=50820 $dt=11
C31 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=40195 $Y=56860 $dt=11
C32 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=40195 $Y=62900 $dt=11
C33 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=40195 $Y=68940 $dt=11
C34 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=41170 $Y=-20340 $dt=11
C35 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=41170 $Y=-8640 $dt=11
C36 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=47210 $Y=-20340 $dt=11
C37 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=47210 $Y=-8640 $dt=11
C38 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=51895 $Y=14580 $dt=11
C39 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=51895 $Y=20620 $dt=11
C40 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=51895 $Y=26660 $dt=11
C41 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=51895 $Y=32700 $dt=11
C42 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=51895 $Y=38740 $dt=11
C43 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=51895 $Y=44780 $dt=11
C44 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=51895 $Y=50820 $dt=11
C45 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=51895 $Y=56860 $dt=11
C46 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=51895 $Y=62900 $dt=11
C47 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=51895 $Y=68940 $dt=11
C48 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=53250 $Y=-20340 $dt=11
C49 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=53250 $Y=-8640 $dt=11
C50 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=59290 $Y=-20340 $dt=11
C51 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=59290 $Y=-8640 $dt=11
C52 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=63595 $Y=14580 $dt=11
C53 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=63595 $Y=20620 $dt=11
C54 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=63595 $Y=26660 $dt=11
C55 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=63595 $Y=32700 $dt=11
C56 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=63595 $Y=38740 $dt=11
C57 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=63595 $Y=44780 $dt=11
C58 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=63595 $Y=50820 $dt=11
C59 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=63595 $Y=56860 $dt=11
C60 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=63595 $Y=62900 $dt=11
C61 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=63595 $Y=68940 $dt=11
C62 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=65330 $Y=-20340 $dt=11
C63 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=65330 $Y=-8640 $dt=11
C64 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=71370 $Y=-20340 $dt=11
C65 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=71370 $Y=-8640 $dt=11
C66 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=75295 $Y=14580 $dt=11
C67 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=75295 $Y=20620 $dt=11
C68 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=75295 $Y=26660 $dt=11
C69 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=75295 $Y=32700 $dt=11
C70 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=75295 $Y=38740 $dt=11
C71 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=75295 $Y=44780 $dt=11
C72 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=75295 $Y=50820 $dt=11
C73 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=75295 $Y=56860 $dt=11
C74 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=75295 $Y=62900 $dt=11
C75 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=75295 $Y=68940 $dt=11
C76 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=77410 $Y=-20340 $dt=11
C77 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=77410 $Y=-8640 $dt=11
C78 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=83450 $Y=-20340 $dt=11
C79 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=83450 $Y=-8640 $dt=11
C80 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=86995 $Y=14580 $dt=11
C81 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=86995 $Y=20620 $dt=11
C82 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=86995 $Y=26660 $dt=11
C83 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=86995 $Y=32700 $dt=11
C84 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=86995 $Y=38740 $dt=11
C85 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=86995 $Y=44780 $dt=11
C86 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=86995 $Y=50820 $dt=11
C87 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=86995 $Y=56860 $dt=11
C88 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=86995 $Y=62900 $dt=11
C89 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=86995 $Y=68940 $dt=11
C90 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=89490 $Y=-20340 $dt=11
C91 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=89490 $Y=-8640 $dt=11
C92 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=95530 $Y=-20340 $dt=11
C93 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=95530 $Y=-8640 $dt=11
C94 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=98695 $Y=14580 $dt=11
C95 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=98695 $Y=20620 $dt=11
C96 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=98695 $Y=26660 $dt=11
C97 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=98695 $Y=32700 $dt=11
C98 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=98695 $Y=38740 $dt=11
C99 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=98695 $Y=44780 $dt=11
C100 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=98695 $Y=50820 $dt=11
C101 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=98695 $Y=56860 $dt=11
C102 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=98695 $Y=62900 $dt=11
C103 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=98695 $Y=68940 $dt=11
C104 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=101570 $Y=-20340 $dt=11
C105 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=101570 $Y=-8640 $dt=11
C106 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=107610 $Y=-20340 $dt=11
C107 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=107610 $Y=-8640 $dt=11
C108 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=110395 $Y=14580 $dt=11
C109 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=110395 $Y=20620 $dt=11
C110 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=110395 $Y=26660 $dt=11
C111 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=110395 $Y=32700 $dt=11
C112 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=110395 $Y=38740 $dt=11
C113 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=110395 $Y=44780 $dt=11
C114 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=110395 $Y=50820 $dt=11
C115 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=110395 $Y=56860 $dt=11
C116 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=110395 $Y=62900 $dt=11
C117 4 3 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=110395 $Y=68940 $dt=11
C118 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=113650 $Y=-20340 $dt=11
C119 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=113650 $Y=-8640 $dt=11
C120 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=119690 $Y=-20340 $dt=11
C121 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=119690 $Y=-8640 $dt=11
C122 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=125730 $Y=-20340 $dt=11
C123 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=125730 $Y=-8640 $dt=11
C124 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=126030 $Y=10220 $dt=11
C125 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=126030 $Y=21920 $dt=11
C126 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=126030 $Y=33620 $dt=11
C127 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=131770 $Y=-20340 $dt=11
C128 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=131770 $Y=-8640 $dt=11
C129 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=132070 $Y=10220 $dt=11
C130 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=132070 $Y=21920 $dt=11
C131 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=132070 $Y=33620 $dt=11
C132 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=137810 $Y=-20340 $dt=11
C133 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=137810 $Y=-8640 $dt=11
C134 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=138110 $Y=10220 $dt=11
C135 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=138110 $Y=21920 $dt=11
C136 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=138110 $Y=33620 $dt=11
C137 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=143850 $Y=-20340 $dt=11
C138 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=143850 $Y=-8640 $dt=11
C139 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=144150 $Y=10220 $dt=11
C140 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=144150 $Y=21920 $dt=11
C141 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=144150 $Y=33620 $dt=11
C142 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=149890 $Y=-20340 $dt=11
C143 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=149890 $Y=-8640 $dt=11
C144 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=150190 $Y=10220 $dt=11
C145 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=150190 $Y=21920 $dt=11
C146 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=150190 $Y=33620 $dt=11
C147 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=155930 $Y=-20340 $dt=11
C148 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=155930 $Y=-8640 $dt=11
C149 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=156230 $Y=10220 $dt=11
C150 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=156230 $Y=21920 $dt=11
C151 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=156230 $Y=33620 $dt=11
C152 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=161970 $Y=-20340 $dt=11
C153 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=161970 $Y=-8640 $dt=11
C154 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=162270 $Y=10220 $dt=11
C155 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=162270 $Y=21920 $dt=11
C156 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=162270 $Y=33620 $dt=11
C157 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=168010 $Y=-20340 $dt=11
C158 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=168010 $Y=-8640 $dt=11
C159 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=168310 $Y=10220 $dt=11
C160 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=168310 $Y=21920 $dt=11
C161 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=168310 $Y=33620 $dt=11
C162 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=174050 $Y=-20340 $dt=11
C163 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=174050 $Y=-8640 $dt=11
C164 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=174350 $Y=10220 $dt=11
C165 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=174350 $Y=21920 $dt=11
C166 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=174350 $Y=33620 $dt=11
C167 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=180090 $Y=-20340 $dt=11
C168 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=180090 $Y=-8640 $dt=11
C169 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=180390 $Y=10220 $dt=11
C170 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=180390 $Y=21920 $dt=11
C171 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=180390 $Y=33620 $dt=11
C172 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=186130 $Y=-20340 $dt=11
C173 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=186130 $Y=-8640 $dt=11
C174 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=186430 $Y=10220 $dt=11
C175 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=186430 $Y=21920 $dt=11
C176 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=186430 $Y=33620 $dt=11
C177 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=192170 $Y=-20340 $dt=11
C178 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=192170 $Y=-8640 $dt=11
C179 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=192470 $Y=10220 $dt=11
C180 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=192470 $Y=21920 $dt=11
C181 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=192470 $Y=33620 $dt=11
C182 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=198210 $Y=-20340 $dt=11
C183 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=198210 $Y=-8640 $dt=11
C184 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=198510 $Y=10220 $dt=11
C185 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=198510 $Y=21920 $dt=11
C186 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=198510 $Y=33620 $dt=11
C187 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=204250 $Y=-20340 $dt=11
C188 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=204250 $Y=-8640 $dt=11
C189 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=204550 $Y=10220 $dt=11
C190 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=204550 $Y=21920 $dt=11
C191 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=204550 $Y=33620 $dt=11
C192 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=210290 $Y=-20340 $dt=11
C193 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=210290 $Y=-8640 $dt=11
C194 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=210590 $Y=10220 $dt=11
C195 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=210590 $Y=21920 $dt=11
C196 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=210590 $Y=33620 $dt=11
C197 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=216330 $Y=-20340 $dt=11
C198 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=216330 $Y=-8640 $dt=11
C199 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=216630 $Y=10220 $dt=11
C200 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=216630 $Y=21920 $dt=11
C201 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=216630 $Y=33620 $dt=11
C202 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=222370 $Y=-20340 $dt=11
C203 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=222370 $Y=-8640 $dt=11
C204 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=222670 $Y=10220 $dt=11
C205 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=222670 $Y=21920 $dt=11
C206 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=222670 $Y=33620 $dt=11
C207 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=228410 $Y=-20340 $dt=11
C208 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=228410 $Y=-8640 $dt=11
C209 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=228710 $Y=10220 $dt=11
C210 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=228710 $Y=21920 $dt=11
C211 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=228710 $Y=33620 $dt=11
C212 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=234450 $Y=-20340 $dt=11
C213 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=234450 $Y=-8640 $dt=11
C214 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=234750 $Y=10220 $dt=11
C215 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=234750 $Y=21920 $dt=11
C216 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=234750 $Y=33620 $dt=11
C217 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=240490 $Y=-20340 $dt=11
C218 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=240490 $Y=-8640 $dt=11
C219 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=240790 $Y=10220 $dt=11
C220 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=240790 $Y=21920 $dt=11
C221 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=240790 $Y=33620 $dt=11
C222 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=246530 $Y=-20340 $dt=11
C223 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=246530 $Y=-8640 $dt=11
C224 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=246830 $Y=10220 $dt=11
C225 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=246830 $Y=21920 $dt=11
C226 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=246830 $Y=33620 $dt=11
C227 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=252570 $Y=-20340 $dt=11
C228 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=252570 $Y=-8640 $dt=11
C229 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=252870 $Y=10220 $dt=11
C230 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=252870 $Y=21920 $dt=11
C231 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=252870 $Y=33620 $dt=11
C232 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=258610 $Y=-20340 $dt=11
C233 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=258610 $Y=-8640 $dt=11
C234 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=258910 $Y=10220 $dt=11
C235 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=258910 $Y=21920 $dt=11
C236 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=258910 $Y=33620 $dt=11
C237 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=264650 $Y=-20340 $dt=11
C238 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=264650 $Y=-8640 $dt=11
C239 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=264950 $Y=10220 $dt=11
C240 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=264950 $Y=21920 $dt=11
C241 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=264950 $Y=33620 $dt=11
C242 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=270690 $Y=-20340 $dt=11
C243 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=270690 $Y=-8640 $dt=11
C244 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=270990 $Y=10220 $dt=11
C245 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=270990 $Y=21920 $dt=11
C246 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=270990 $Y=33620 $dt=11
C247 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=276730 $Y=-20340 $dt=11
C248 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=276730 $Y=-8640 $dt=11
C249 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=277030 $Y=10220 $dt=11
C250 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=277030 $Y=21920 $dt=11
C251 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=277030 $Y=33620 $dt=11
C252 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=282770 $Y=-20340 $dt=11
C253 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=282770 $Y=-8640 $dt=11
C254 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=283070 $Y=10220 $dt=11
C255 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=283070 $Y=21920 $dt=11
C256 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=283070 $Y=33620 $dt=11
C257 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=288810 $Y=-20340 $dt=11
C258 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=288810 $Y=-8640 $dt=11
C259 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=289110 $Y=10220 $dt=11
C260 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=289110 $Y=21920 $dt=11
C261 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=289110 $Y=33620 $dt=11
C262 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=294850 $Y=-20340 $dt=11
C263 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=294850 $Y=-8640 $dt=11
C264 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=295150 $Y=10220 $dt=11
C265 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=295150 $Y=21920 $dt=11
C266 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=295150 $Y=33620 $dt=11
C267 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=300890 $Y=-20340 $dt=11
C268 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=300890 $Y=-8640 $dt=11
C269 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=301190 $Y=10220 $dt=11
C270 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=301190 $Y=21920 $dt=11
C271 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=301190 $Y=33620 $dt=11
C272 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=306930 $Y=-20340 $dt=11
C273 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=306930 $Y=-8640 $dt=11
C274 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=307230 $Y=10220 $dt=11
C275 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=307230 $Y=21920 $dt=11
C276 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=307230 $Y=33620 $dt=11
C277 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=312970 $Y=-20340 $dt=11
C278 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=312970 $Y=-8640 $dt=11
C279 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=313270 $Y=10220 $dt=11
C280 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=313270 $Y=21920 $dt=11
C281 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=313270 $Y=33620 $dt=11
C282 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=319010 $Y=-20340 $dt=11
C283 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=319010 $Y=-8640 $dt=11
C284 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=319310 $Y=10220 $dt=11
C285 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=319310 $Y=21920 $dt=11
C286 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=319310 $Y=33620 $dt=11
C287 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=325050 $Y=-20340 $dt=11
C288 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=325050 $Y=-8640 $dt=11
C289 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=325350 $Y=10220 $dt=11
C290 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=325350 $Y=21920 $dt=11
C291 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=325350 $Y=33620 $dt=11
C292 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=331090 $Y=-20340 $dt=11
C293 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=331090 $Y=-8640 $dt=11
C294 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=331390 $Y=10220 $dt=11
C295 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=331390 $Y=21920 $dt=11
C296 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=331390 $Y=33620 $dt=11
C297 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=337130 $Y=-20340 $dt=11
C298 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=337130 $Y=-8640 $dt=11
C299 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=337430 $Y=10220 $dt=11
C300 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=337430 $Y=21920 $dt=11
C301 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=337430 $Y=33620 $dt=11
C302 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=343170 $Y=-20340 $dt=11
C303 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=343170 $Y=-8640 $dt=11
C304 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=343470 $Y=10220 $dt=11
C305 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=343470 $Y=21920 $dt=11
C306 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=343470 $Y=33620 $dt=11
C307 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=349210 $Y=-20340 $dt=11
C308 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=349210 $Y=-8640 $dt=11
C309 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=349510 $Y=10220 $dt=11
C310 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=349510 $Y=21920 $dt=11
C311 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=349510 $Y=33620 $dt=11
C312 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=355250 $Y=-20340 $dt=11
C313 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=355250 $Y=-8640 $dt=11
C314 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=355550 $Y=10220 $dt=11
C315 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=355550 $Y=21920 $dt=11
C316 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=355550 $Y=33620 $dt=11
C317 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=361290 $Y=-20340 $dt=11
C318 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=361290 $Y=-8640 $dt=11
C319 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=361590 $Y=10220 $dt=11
C320 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=361590 $Y=21920 $dt=11
C321 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=361590 $Y=33620 $dt=11
C322 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=367330 $Y=-20340 $dt=11
C323 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=367330 $Y=-8640 $dt=11
C324 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=367630 $Y=10220 $dt=11
C325 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=367630 $Y=21920 $dt=11
C326 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=367630 $Y=33620 $dt=11
C327 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=373370 $Y=-20340 $dt=11
C328 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=373370 $Y=-8640 $dt=11
C329 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=373670 $Y=10220 $dt=11
C330 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=373670 $Y=21920 $dt=11
C331 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=373670 $Y=33620 $dt=11
C332 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=379410 $Y=-20340 $dt=11
C333 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=379410 $Y=-8640 $dt=11
C334 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=379710 $Y=10220 $dt=11
C335 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=379710 $Y=21920 $dt=11
C336 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=379710 $Y=33620 $dt=11
C337 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=385450 $Y=-20340 $dt=11
C338 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=385450 $Y=-8640 $dt=11
C339 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=385750 $Y=10220 $dt=11
C340 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=385750 $Y=21920 $dt=11
C341 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=385750 $Y=33620 $dt=11
C342 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=391490 $Y=-20340 $dt=11
C343 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=391490 $Y=-8640 $dt=11
C344 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=391790 $Y=10220 $dt=11
C345 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=391790 $Y=21920 $dt=11
C346 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=391790 $Y=33620 $dt=11
C347 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=397530 $Y=-20340 $dt=11
C348 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=397530 $Y=-8640 $dt=11
C349 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=397830 $Y=10220 $dt=11
C350 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=397830 $Y=21920 $dt=11
C351 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=397830 $Y=33620 $dt=11
C352 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=403570 $Y=-20340 $dt=11
C353 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=403570 $Y=-8640 $dt=11
C354 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=403870 $Y=10220 $dt=11
C355 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=403870 $Y=21920 $dt=11
C356 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=403870 $Y=33620 $dt=11
C357 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=409610 $Y=-20340 $dt=11
C358 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=409610 $Y=-8640 $dt=11
C359 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=409910 $Y=10220 $dt=11
C360 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=409910 $Y=21920 $dt=11
C361 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=409910 $Y=33620 $dt=11
C362 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=415650 $Y=-20340 $dt=11
C363 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=415650 $Y=-8640 $dt=11
C364 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=415950 $Y=10220 $dt=11
C365 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=415950 $Y=21920 $dt=11
C366 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=415950 $Y=33620 $dt=11
C367 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=421690 $Y=-20340 $dt=11
C368 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=421690 $Y=-8640 $dt=11
C369 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=421990 $Y=10220 $dt=11
C370 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=421990 $Y=21920 $dt=11
C371 2 1 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=421990 $Y=33620 $dt=11
.ends MASCO__P4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_723062655414                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_723062655414 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_723062655414

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_723062655418                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_723062655418 1 2
** N=2 EP=2 FDC=0
.ends VIA1_C_CDNS_723062655418

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_723062655419                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_723062655419 1 2
** N=2 EP=2 FDC=0
.ends VIA1_C_CDNS_723062655419

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7230626554120                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7230626554120 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7230626554120

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_7230626554124                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_7230626554124 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_7230626554124

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_7230626554125                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_7230626554125 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_7230626554125

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7230626554127                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7230626554127 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7230626554127

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_7230626554128                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_7230626554128 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_7230626554128

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_7230626554129                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_7230626554129 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_7230626554129

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_7230626554130                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_7230626554130 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_7230626554130

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_7230626554132                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_7230626554132 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_7230626554132

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_7230626554133                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_7230626554133 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_7230626554133

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7230626554138                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7230626554138 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7230626554138

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7230626554139                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7230626554139 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7230626554139

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7230626554140                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7230626554140 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7230626554140

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7230626554142                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7230626554142 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7230626554142

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7230626554144                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7230626554144 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7230626554144

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7230626554147                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7230626554147 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7230626554147

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ped_CDNS_723062655411                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ped_CDNS_723062655411 1 2 3 4
** N=4 EP=4 FDC=12
X0 2 4 3 1 LDDP w=5e-05 l=9.4e-07 ad=2.19714e-10 pd=8.94366e-05 adio=4.2498e-10 pdio=2.57015e-05 extlay=1 $[ped] $X=-2270 $Y=0 $dt=1
X1 2 4 3 1 LDDP w=5e-05 l=9.4e-07 ad=2.19714e-10 pd=8.94366e-05 adio=4.2498e-10 pdio=2.57015e-05 extlay=1 $[ped] $X=6530 $Y=0 $dt=1
X2 2 4 3 1 LDDP w=5e-05 l=9.4e-07 ad=2.19714e-10 pd=8.94366e-05 adio=4.2498e-10 pdio=2.57015e-05 extlay=1 $[ped] $X=15330 $Y=0 $dt=1
X3 2 4 3 1 LDDP w=5e-05 l=9.4e-07 ad=2.19714e-10 pd=8.94366e-05 adio=4.2498e-10 pdio=2.57015e-05 extlay=1 $[ped] $X=24130 $Y=0 $dt=1
X4 2 4 3 1 LDDP w=5e-05 l=9.4e-07 ad=2.19714e-10 pd=8.94366e-05 adio=4.2498e-10 pdio=2.57015e-05 extlay=1 $[ped] $X=32930 $Y=0 $dt=1
X5 2 4 3 1 LDDP w=5e-05 l=9.4e-07 ad=2.19714e-10 pd=8.94366e-05 adio=4.2498e-10 pdio=2.57015e-05 extlay=1 $[ped] $X=41730 $Y=0 $dt=1
X6 2 4 3 1 LDDP w=5e-05 l=9.4e-07 ad=2.19714e-10 pd=8.94366e-05 adio=4.2498e-10 pdio=2.57015e-05 extlay=1 $[ped] $X=50530 $Y=0 $dt=1
X7 2 4 3 1 LDDP w=5e-05 l=9.4e-07 ad=2.19714e-10 pd=8.94366e-05 adio=4.2498e-10 pdio=2.57015e-05 extlay=1 $[ped] $X=59330 $Y=0 $dt=1
X8 2 4 3 1 LDDP w=5e-05 l=9.4e-07 ad=2.19714e-10 pd=8.94366e-05 adio=4.2498e-10 pdio=2.57015e-05 extlay=1 $[ped] $X=68130 $Y=0 $dt=1
X9 2 4 3 1 LDDP w=5e-05 l=9.4e-07 ad=2.19714e-10 pd=8.94366e-05 adio=4.2498e-10 pdio=2.57015e-05 extlay=1 $[ped] $X=76930 $Y=0 $dt=1
X10 2 4 3 1 LDDP w=5e-05 l=9.4e-07 ad=2.19714e-10 pd=8.94366e-05 adio=4.2498e-10 pdio=2.57015e-05 extlay=1 $[ped] $X=85730 $Y=0 $dt=1
X11 2 4 3 1 LDDP w=5e-05 l=9.4e-07 ad=2.19714e-10 pd=8.94366e-05 adio=4.2498e-10 pdio=2.57015e-05 extlay=1 $[ped] $X=94530 $Y=0 $dt=1
.ends ped_CDNS_723062655411

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_723062655412                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_723062655412 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.00204358 W=2e-06 $[rpp1k1_3] $SUB=3 $X=-2220 $Y=0 $dt=10
.ends rpp1k1_3_CDNS_723062655412

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_723062655416                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_723062655416 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.0002029 W=2e-06 $[rpp1k1_3] $SUB=3 $X=-2220 $Y=0 $dt=10
.ends rpp1k1_3_CDNS_723062655416

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: dpp20_CDNS_723062655418                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt dpp20_CDNS_723062655418 1 2 3
** N=3 EP=3 FDC=2
D0 1 2 p_ddnw AREA=1.12107e-09 PJ=0.00016136 perimeter=0.00016136 $X=-6420 $Y=-6420 $dt=5
D1 3 2 dpp20 AREA=2.5e-10 PJ=0.00011 perimeter=0.00011 $X=0 $Y=0 $dt=7
.ends dpp20_CDNS_723062655418

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_723062655419                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_723062655419 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.0002537 W=2e-06 $[rpp1k1_3] $SUB=3 $X=-2220 $Y=0 $dt=10
.ends rpp1k1_3_CDNS_723062655419

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X13                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X13 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7230626554116 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7230626554116 $T=500 1500 0 0 $X=0 $Y=1000
X2 1 VIATP_C_CDNS_7230626554116 $T=500 2500 0 0 $X=0 $Y=2000
X3 1 VIATP_C_CDNS_7230626554116 $T=500 3500 0 0 $X=0 $Y=3000
X4 1 VIATP_C_CDNS_7230626554116 $T=500 4500 0 0 $X=0 $Y=4000
X5 1 VIATP_C_CDNS_7230626554116 $T=500 5500 0 0 $X=0 $Y=5000
X6 1 VIATP_C_CDNS_7230626554116 $T=500 6500 0 0 $X=0 $Y=6000
.ends MASCO__X13

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y15                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y15 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7230626554140 $T=500 440 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7230626554140 $T=1500 440 0 0 $X=1000 $Y=0
X2 1 VIATP_C_CDNS_7230626554140 $T=2500 440 0 0 $X=2000 $Y=0
X3 1 VIATP_C_CDNS_7230626554140 $T=3500 440 0 0 $X=3000 $Y=0
X4 1 VIATP_C_CDNS_7230626554140 $T=4500 440 0 0 $X=4000 $Y=0
X5 1 VIATP_C_CDNS_7230626554140 $T=5500 440 0 0 $X=5000 $Y=0
X6 1 VIATP_C_CDNS_7230626554140 $T=6500 440 0 0 $X=6000 $Y=0
X7 1 VIATP_C_CDNS_7230626554140 $T=7500 440 0 0 $X=7000 $Y=0
X8 1 VIATP_C_CDNS_7230626554140 $T=8500 440 0 0 $X=8000 $Y=0
X9 1 VIATP_C_CDNS_7230626554140 $T=9500 440 0 0 $X=9000 $Y=0
X10 1 VIATP_C_CDNS_7230626554140 $T=10500 440 0 0 $X=10000 $Y=0
X11 1 VIATP_C_CDNS_7230626554140 $T=11500 440 0 0 $X=11000 $Y=0
.ends MASCO__Y15

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X11                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X11 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7230626554116 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7230626554116 $T=500 2500 0 0 $X=0 $Y=2000
X2 1 VIATP_C_CDNS_7230626554116 $T=500 4500 0 0 $X=0 $Y=4000
X3 1 VIATP_C_CDNS_7230626554116 $T=500 6500 0 0 $X=0 $Y=6000
X4 1 VIATP_C_CDNS_7230626554116 $T=500 8500 0 0 $X=0 $Y=8000
X5 1 VIATP_C_CDNS_7230626554116 $T=500 10500 0 0 $X=0 $Y=10000
X6 1 VIATP_C_CDNS_7230626554116 $T=500 12500 0 0 $X=0 $Y=12000
X7 1 VIATP_C_CDNS_7230626554116 $T=500 14500 0 0 $X=0 $Y=14000
X8 1 VIATP_C_CDNS_7230626554116 $T=500 16500 0 0 $X=0 $Y=16000
.ends MASCO__X11

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y16                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y16 1
** N=1 EP=1 FDC=0
X0 1 MASCO__X11 $T=0 0 0 0 $X=0 $Y=0
X1 1 MASCO__X11 $T=2000 0 0 0 $X=2000 $Y=0
X2 1 MASCO__X11 $T=4000 0 0 0 $X=4000 $Y=0
X3 1 MASCO__X11 $T=6000 0 0 0 $X=6000 $Y=0
.ends MASCO__Y16

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y17                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y17 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7230626554136 $T=500 620 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7230626554136 $T=1500 620 0 0 $X=1000 $Y=0
X2 1 VIATP_C_CDNS_7230626554136 $T=2500 620 0 0 $X=2000 $Y=0
X3 1 VIATP_C_CDNS_7230626554136 $T=3500 620 0 0 $X=3000 $Y=0
X4 1 VIATP_C_CDNS_7230626554136 $T=4500 620 0 0 $X=4000 $Y=0
X5 1 VIATP_C_CDNS_7230626554136 $T=5500 620 0 0 $X=5000 $Y=0
.ends MASCO__Y17

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y19                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y19 1
** N=1 EP=1 FDC=0
X0 1 MASCO__X8 $T=0 0 0 0 $X=0 $Y=0
X1 1 MASCO__X8 $T=2000 0 0 0 $X=2000 $Y=0
X2 1 MASCO__X8 $T=4000 0 0 0 $X=4000 $Y=0
X3 1 MASCO__X8 $T=6000 0 0 0 $X=6000 $Y=0
.ends MASCO__Y19

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y20                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y20 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7230626554134 $T=500 750 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7230626554134 $T=1500 750 0 0 $X=1000 $Y=0
X2 1 VIATP_C_CDNS_7230626554134 $T=2500 750 0 0 $X=2000 $Y=0
X3 1 VIATP_C_CDNS_7230626554134 $T=3500 750 0 0 $X=3000 $Y=0
X4 1 VIATP_C_CDNS_7230626554134 $T=4500 750 0 0 $X=4000 $Y=0
X5 1 VIATP_C_CDNS_7230626554134 $T=5500 750 0 0 $X=5000 $Y=0
X6 1 VIATP_C_CDNS_7230626554134 $T=6500 750 0 0 $X=6000 $Y=0
X7 1 VIATP_C_CDNS_7230626554134 $T=7500 750 0 0 $X=7000 $Y=0
.ends MASCO__Y20

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y21                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y21 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7230626554116 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7230626554116 $T=2500 500 0 0 $X=2000 $Y=0
X2 1 VIATP_C_CDNS_7230626554116 $T=4500 500 0 0 $X=4000 $Y=0
X3 1 VIATP_C_CDNS_7230626554116 $T=6500 500 0 0 $X=6000 $Y=0
.ends MASCO__Y21

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__P5                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__P5 1 2 3 4 5 6
** N=7 EP=6 FDC=21
X0 1 VIA1_C_CDNS_723062655414 $T=42315 186985 0 0 $X=41565 $Y=185975
X1 2 VIA1_C_CDNS_723062655414 $T=46630 168085 0 0 $X=45880 $Y=167075
X2 3 VIA1_C_CDNS_723062655414 $T=48475 149805 0 0 $X=47725 $Y=148795
X3 4 VIA1_C_CDNS_723062655414 $T=82400 149805 0 0 $X=81650 $Y=148795
X4 1 VIA1_C_CDNS_723062655414 $T=88760 186595 0 0 $X=88010 $Y=185585
X5 1 6 VIA1_C_CDNS_723062655418 $T=168435 182510 0 0 $X=158065 $Y=182020
X6 1 6 VIA1_C_CDNS_723062655418 $T=245255 182765 0 0 $X=234885 $Y=182275
X7 5 6 VIA1_C_CDNS_723062655419 $T=167770 176605 0 0 $X=143240 $Y=174710
X8 5 6 VIA1_C_CDNS_723062655419 $T=245135 176605 0 0 $X=220605 $Y=174710
X9 1 VIATP_C_CDNS_7230626554120 $T=298975 183945 0 0 $X=298100 $Y=183445
X10 1 VIATP_C_CDNS_7230626554120 $T=298975 184945 0 0 $X=298100 $Y=184445
X11 1 VIATP_C_CDNS_7230626554120 $T=298975 185945 0 0 $X=298100 $Y=185445
X12 1 VIATP_C_CDNS_7230626554120 $T=298975 186945 0 0 $X=298100 $Y=186445
X13 1 VIATP_C_CDNS_7230626554120 $T=298975 187945 0 0 $X=298100 $Y=187445
X14 1 VIATP_C_CDNS_7230626554120 $T=298975 188945 0 0 $X=298100 $Y=188445
X15 1 VIATP_C_CDNS_7230626554120 $T=298975 189945 0 0 $X=298100 $Y=189445
X16 1 VIATP_C_CDNS_7230626554120 $T=298975 191945 0 0 $X=298100 $Y=191445
X17 1 VIATP_C_CDNS_7230626554120 $T=298975 192945 0 0 $X=298100 $Y=192445
X18 1 VIATP_C_CDNS_7230626554120 $T=298975 193945 0 0 $X=298100 $Y=193445
X19 1 VIATP_C_CDNS_7230626554120 $T=298975 194945 0 0 $X=298100 $Y=194445
X20 1 VIATP_C_CDNS_7230626554120 $T=298975 195945 0 0 $X=298100 $Y=195445
X21 1 VIATP_C_CDNS_7230626554120 $T=298975 196945 0 0 $X=298100 $Y=196445
X22 1 VIATP_C_CDNS_7230626554120 $T=298975 197945 0 0 $X=298100 $Y=197445
X23 1 VIATP_C_CDNS_7230626554120 $T=298975 198945 0 0 $X=298100 $Y=198445
X24 1 VIATP_C_CDNS_7230626554120 $T=298975 199945 0 0 $X=298100 $Y=199445
X25 1 VIATP_C_CDNS_7230626554120 $T=298975 200945 0 0 $X=298100 $Y=200445
X26 1 VIATP_C_CDNS_7230626554120 $T=298975 201945 0 0 $X=298100 $Y=201445
X27 1 VIATP_C_CDNS_7230626554120 $T=298975 202945 0 0 $X=298100 $Y=202445
X28 1 VIATP_C_CDNS_7230626554120 $T=298975 203945 0 0 $X=298100 $Y=203445
X29 1 VIATP_C_CDNS_7230626554120 $T=298975 204945 0 0 $X=298100 $Y=204445
X30 1 VIATP_C_CDNS_7230626554120 $T=298975 206945 0 0 $X=298100 $Y=206445
X31 1 VIATP_C_CDNS_7230626554120 $T=298975 207945 0 0 $X=298100 $Y=207445
X32 1 VIATP_C_CDNS_7230626554120 $T=298975 208945 0 0 $X=298100 $Y=208445
X33 1 VIATP_C_CDNS_7230626554120 $T=298975 209945 0 0 $X=298100 $Y=209445
X34 1 VIATP_C_CDNS_7230626554120 $T=433725 183945 0 0 $X=432850 $Y=183445
X35 1 VIATP_C_CDNS_7230626554120 $T=433725 184945 0 0 $X=432850 $Y=184445
X36 1 VIATP_C_CDNS_7230626554120 $T=433725 185945 0 0 $X=432850 $Y=185445
X37 1 VIATP_C_CDNS_7230626554120 $T=433725 186945 0 0 $X=432850 $Y=186445
X38 1 VIATP_C_CDNS_7230626554120 $T=433725 187945 0 0 $X=432850 $Y=187445
X39 1 VIATP_C_CDNS_7230626554120 $T=433725 188945 0 0 $X=432850 $Y=188445
X40 1 VIATP_C_CDNS_7230626554120 $T=433725 189945 0 0 $X=432850 $Y=189445
X41 1 VIATP_C_CDNS_7230626554120 $T=433725 190945 0 0 $X=432850 $Y=190445
X42 1 VIATP_C_CDNS_7230626554120 $T=433725 191945 0 0 $X=432850 $Y=191445
X43 1 VIATP_C_CDNS_7230626554120 $T=433725 192945 0 0 $X=432850 $Y=192445
X44 1 VIATP_C_CDNS_7230626554120 $T=433725 193945 0 0 $X=432850 $Y=193445
X45 1 VIATP_C_CDNS_7230626554120 $T=433725 194945 0 0 $X=432850 $Y=194445
X46 1 VIATP_C_CDNS_7230626554120 $T=433725 195945 0 0 $X=432850 $Y=195445
X47 1 VIATP_C_CDNS_7230626554120 $T=433725 196945 0 0 $X=432850 $Y=196445
X48 1 VIATP_C_CDNS_7230626554120 $T=433725 197945 0 0 $X=432850 $Y=197445
X49 1 VIATP_C_CDNS_7230626554120 $T=433725 198945 0 0 $X=432850 $Y=198445
X50 1 VIATP_C_CDNS_7230626554120 $T=433725 199945 0 0 $X=432850 $Y=199445
X51 1 VIATP_C_CDNS_7230626554120 $T=433725 200945 0 0 $X=432850 $Y=200445
X52 1 VIATP_C_CDNS_7230626554120 $T=433725 201945 0 0 $X=432850 $Y=201445
X53 1 VIATP_C_CDNS_7230626554120 $T=433725 202945 0 0 $X=432850 $Y=202445
X54 1 VIATP_C_CDNS_7230626554120 $T=433725 203945 0 0 $X=432850 $Y=203445
X55 1 VIATP_C_CDNS_7230626554120 $T=433725 204945 0 0 $X=432850 $Y=204445
X56 1 VIATP_C_CDNS_7230626554120 $T=433725 205945 0 0 $X=432850 $Y=205445
X57 1 VIATP_C_CDNS_7230626554120 $T=433725 206945 0 0 $X=432850 $Y=206445
X58 1 VIATP_C_CDNS_7230626554120 $T=433725 207945 0 0 $X=432850 $Y=207445
X59 1 VIATP_C_CDNS_7230626554120 $T=433725 208945 0 0 $X=432850 $Y=208445
X60 1 VIATP_C_CDNS_7230626554120 $T=433725 209945 0 0 $X=432850 $Y=209445
X61 5 VIA3_C_CDNS_7230626554124 $T=261795 138745 0 0 $X=261060 $Y=138245
X62 5 VIA3_C_CDNS_7230626554124 $T=261795 140745 0 0 $X=261060 $Y=140245
X63 5 VIA3_C_CDNS_7230626554124 $T=261795 142745 0 0 $X=261060 $Y=142245
X64 5 VIA3_C_CDNS_7230626554124 $T=261795 144745 0 0 $X=261060 $Y=144245
X65 5 VIA3_C_CDNS_7230626554125 $T=264035 137745 0 0 $X=263535 $Y=137245
X66 5 VIA3_C_CDNS_7230626554125 $T=264035 139745 0 0 $X=263535 $Y=139245
X67 5 VIA3_C_CDNS_7230626554125 $T=264035 141745 0 0 $X=263535 $Y=141245
X68 5 VIA3_C_CDNS_7230626554125 $T=264035 143745 0 0 $X=263535 $Y=143245
X69 5 VIA3_C_CDNS_7230626554125 $T=266035 137745 0 0 $X=265535 $Y=137245
X70 5 VIA3_C_CDNS_7230626554125 $T=266035 139745 0 0 $X=265535 $Y=139245
X71 5 VIA3_C_CDNS_7230626554125 $T=266035 141745 0 0 $X=265535 $Y=141245
X72 5 VIA3_C_CDNS_7230626554125 $T=266035 143745 0 0 $X=265535 $Y=143245
X73 5 VIA3_C_CDNS_7230626554125 $T=268035 137745 0 0 $X=267535 $Y=137245
X74 5 VIA3_C_CDNS_7230626554125 $T=268035 139745 0 0 $X=267535 $Y=139245
X75 5 VIA3_C_CDNS_7230626554125 $T=268035 141745 0 0 $X=267535 $Y=141245
X76 5 VIA3_C_CDNS_7230626554125 $T=268035 143745 0 0 $X=267535 $Y=143245
X77 5 VIA3_C_CDNS_7230626554125 $T=270035 137745 0 0 $X=269535 $Y=137245
X78 5 VIA3_C_CDNS_7230626554125 $T=270035 139745 0 0 $X=269535 $Y=139245
X79 5 VIA3_C_CDNS_7230626554125 $T=270035 141745 0 0 $X=269535 $Y=141245
X80 5 VIA3_C_CDNS_7230626554125 $T=270035 143745 0 0 $X=269535 $Y=143245
X81 1 VIATP_C_CDNS_7230626554127 $T=405105 183945 0 0 $X=404835 $Y=183445
X82 1 VIATP_C_CDNS_7230626554127 $T=405105 184945 0 0 $X=404835 $Y=184445
X83 1 VIATP_C_CDNS_7230626554127 $T=405105 185945 0 0 $X=404835 $Y=185445
X84 1 VIATP_C_CDNS_7230626554127 $T=405105 186945 0 0 $X=404835 $Y=186445
X85 1 VIATP_C_CDNS_7230626554127 $T=405105 187945 0 0 $X=404835 $Y=187445
X86 1 VIATP_C_CDNS_7230626554127 $T=405105 188945 0 0 $X=404835 $Y=188445
X87 1 VIATP_C_CDNS_7230626554127 $T=405105 189945 0 0 $X=404835 $Y=189445
X88 1 VIATP_C_CDNS_7230626554127 $T=405105 190945 0 0 $X=404835 $Y=190445
X89 1 VIATP_C_CDNS_7230626554127 $T=405105 191945 0 0 $X=404835 $Y=191445
X90 1 VIATP_C_CDNS_7230626554127 $T=405105 192945 0 0 $X=404835 $Y=192445
X91 1 VIATP_C_CDNS_7230626554127 $T=405105 193945 0 0 $X=404835 $Y=193445
X92 1 VIATP_C_CDNS_7230626554127 $T=405105 194945 0 0 $X=404835 $Y=194445
X93 1 VIATP_C_CDNS_7230626554127 $T=405105 195945 0 0 $X=404835 $Y=195445
X94 1 VIATP_C_CDNS_7230626554127 $T=405105 196945 0 0 $X=404835 $Y=196445
X95 1 VIATP_C_CDNS_7230626554127 $T=405105 197945 0 0 $X=404835 $Y=197445
X96 1 VIATP_C_CDNS_7230626554127 $T=405105 198945 0 0 $X=404835 $Y=198445
X97 1 VIATP_C_CDNS_7230626554127 $T=405105 199945 0 0 $X=404835 $Y=199445
X98 1 VIATP_C_CDNS_7230626554127 $T=405105 200945 0 0 $X=404835 $Y=200445
X99 1 VIATP_C_CDNS_7230626554127 $T=405105 201945 0 0 $X=404835 $Y=201445
X100 1 VIATP_C_CDNS_7230626554127 $T=405105 202945 0 0 $X=404835 $Y=202445
X101 1 VIATP_C_CDNS_7230626554127 $T=405105 203945 0 0 $X=404835 $Y=203445
X102 1 VIATP_C_CDNS_7230626554127 $T=405105 204945 0 0 $X=404835 $Y=204445
X103 1 VIATP_C_CDNS_7230626554127 $T=405105 205945 0 0 $X=404835 $Y=205445
X104 1 VIATP_C_CDNS_7230626554127 $T=405105 206945 0 0 $X=404835 $Y=206445
X105 1 VIATP_C_CDNS_7230626554127 $T=405105 207945 0 0 $X=404835 $Y=207445
X106 1 VIATP_C_CDNS_7230626554127 $T=405105 208945 0 0 $X=404835 $Y=208445
X107 1 VIATP_C_CDNS_7230626554127 $T=405105 209945 0 0 $X=404835 $Y=209445
X108 5 VIA3_C_CDNS_7230626554128 $T=261795 137745 0 0 $X=261060 $Y=137245
X109 5 VIA3_C_CDNS_7230626554128 $T=261795 139745 0 0 $X=261060 $Y=139245
X110 5 VIA3_C_CDNS_7230626554128 $T=261795 141745 0 0 $X=261060 $Y=141245
X111 5 VIA3_C_CDNS_7230626554128 $T=261795 143745 0 0 $X=261060 $Y=143245
X112 5 VIA3_C_CDNS_7230626554129 $T=263035 137745 0 0 $X=262535 $Y=137245
X113 5 VIA3_C_CDNS_7230626554129 $T=263035 139745 0 0 $X=262535 $Y=139245
X114 5 VIA3_C_CDNS_7230626554129 $T=263035 141745 0 0 $X=262535 $Y=141245
X115 5 VIA3_C_CDNS_7230626554129 $T=263035 143745 0 0 $X=262535 $Y=143245
X116 5 VIA3_C_CDNS_7230626554129 $T=265035 137745 0 0 $X=264535 $Y=137245
X117 5 VIA3_C_CDNS_7230626554129 $T=265035 139745 0 0 $X=264535 $Y=139245
X118 5 VIA3_C_CDNS_7230626554129 $T=265035 141745 0 0 $X=264535 $Y=141245
X119 5 VIA3_C_CDNS_7230626554129 $T=265035 143745 0 0 $X=264535 $Y=143245
X120 5 VIA3_C_CDNS_7230626554129 $T=267035 137745 0 0 $X=266535 $Y=137245
X121 5 VIA3_C_CDNS_7230626554129 $T=267035 139745 0 0 $X=266535 $Y=139245
X122 5 VIA3_C_CDNS_7230626554129 $T=267035 141745 0 0 $X=266535 $Y=141245
X123 5 VIA3_C_CDNS_7230626554129 $T=267035 143745 0 0 $X=266535 $Y=143245
X124 5 VIA3_C_CDNS_7230626554129 $T=269035 137745 0 0 $X=268535 $Y=137245
X125 5 VIA3_C_CDNS_7230626554129 $T=269035 139745 0 0 $X=268535 $Y=139245
X126 5 VIA3_C_CDNS_7230626554129 $T=269035 141745 0 0 $X=268535 $Y=141245
X127 5 VIA3_C_CDNS_7230626554129 $T=269035 143745 0 0 $X=268535 $Y=143245
X128 5 VIA3_C_CDNS_7230626554130 $T=264035 138745 0 0 $X=263535 $Y=138245
X129 5 VIA3_C_CDNS_7230626554130 $T=264035 140745 0 0 $X=263535 $Y=140245
X130 5 VIA3_C_CDNS_7230626554130 $T=264035 142745 0 0 $X=263535 $Y=142245
X131 5 VIA3_C_CDNS_7230626554130 $T=264035 144745 0 0 $X=263535 $Y=144245
X132 5 VIA3_C_CDNS_7230626554130 $T=266035 138745 0 0 $X=265535 $Y=138245
X133 5 VIA3_C_CDNS_7230626554130 $T=266035 140745 0 0 $X=265535 $Y=140245
X134 5 VIA3_C_CDNS_7230626554130 $T=266035 142745 0 0 $X=265535 $Y=142245
X135 5 VIA3_C_CDNS_7230626554130 $T=266035 144745 0 0 $X=265535 $Y=144245
X136 5 VIA3_C_CDNS_7230626554130 $T=268035 138745 0 0 $X=267535 $Y=138245
X137 5 VIA3_C_CDNS_7230626554130 $T=268035 140745 0 0 $X=267535 $Y=140245
X138 5 VIA3_C_CDNS_7230626554130 $T=268035 142745 0 0 $X=267535 $Y=142245
X139 5 VIA3_C_CDNS_7230626554130 $T=268035 144745 0 0 $X=267535 $Y=144245
X140 5 VIA3_C_CDNS_7230626554130 $T=270035 138745 0 0 $X=269535 $Y=138245
X141 5 VIA3_C_CDNS_7230626554130 $T=270035 140745 0 0 $X=269535 $Y=140245
X142 5 VIA3_C_CDNS_7230626554130 $T=270035 142745 0 0 $X=269535 $Y=142245
X143 5 VIA3_C_CDNS_7230626554130 $T=270035 144745 0 0 $X=269535 $Y=144245
X144 5 VIA3_C_CDNS_7230626554132 $T=263035 145995 0 0 $X=262535 $Y=145245
X145 5 VIA3_C_CDNS_7230626554132 $T=265035 145995 0 0 $X=264535 $Y=145245
X146 5 VIA3_C_CDNS_7230626554132 $T=267035 145995 0 0 $X=266535 $Y=145245
X147 5 VIA3_C_CDNS_7230626554132 $T=269035 145995 0 0 $X=268535 $Y=145245
X148 5 VIA3_C_CDNS_7230626554133 $T=264035 145995 0 0 $X=263535 $Y=145245
X149 5 VIA3_C_CDNS_7230626554133 $T=266035 145995 0 0 $X=265535 $Y=145245
X150 5 VIA3_C_CDNS_7230626554133 $T=268035 145995 0 0 $X=267535 $Y=145245
X151 5 VIA3_C_CDNS_7230626554133 $T=270035 145995 0 0 $X=269535 $Y=145245
X152 1 VIATP_C_CDNS_7230626554134 $T=406350 211195 0 0 $X=405850 $Y=210445
X153 1 VIATP_C_CDNS_7230626554134 $T=407350 211195 0 0 $X=406850 $Y=210445
X154 1 VIATP_C_CDNS_7230626554134 $T=408350 211195 0 0 $X=407850 $Y=210445
X155 1 VIATP_C_CDNS_7230626554134 $T=409350 211195 0 0 $X=408850 $Y=210445
X156 1 VIATP_C_CDNS_7230626554134 $T=410350 211195 0 0 $X=409850 $Y=210445
X157 1 VIATP_C_CDNS_7230626554134 $T=411350 211195 0 0 $X=410850 $Y=210445
X158 1 VIATP_C_CDNS_7230626554134 $T=412350 211195 0 0 $X=411850 $Y=210445
X159 1 VIATP_C_CDNS_7230626554134 $T=413350 211195 0 0 $X=412850 $Y=210445
X160 1 VIATP_C_CDNS_7230626554134 $T=414350 211195 0 0 $X=413850 $Y=210445
X161 1 VIATP_C_CDNS_7230626554134 $T=415350 211195 0 0 $X=414850 $Y=210445
X162 1 VIATP_C_CDNS_7230626554134 $T=416350 211195 0 0 $X=415850 $Y=210445
X163 1 VIATP_C_CDNS_7230626554134 $T=417350 211195 0 0 $X=416850 $Y=210445
X164 1 VIATP_C_CDNS_7230626554134 $T=418350 211195 0 0 $X=417850 $Y=210445
X165 1 VIATP_C_CDNS_7230626554134 $T=419350 211195 0 0 $X=418850 $Y=210445
X166 1 VIATP_C_CDNS_7230626554134 $T=420350 211195 0 0 $X=419850 $Y=210445
X167 1 VIATP_C_CDNS_7230626554134 $T=421350 211195 0 0 $X=420850 $Y=210445
X168 1 VIATP_C_CDNS_7230626554134 $T=422350 211195 0 0 $X=421850 $Y=210445
X169 1 VIATP_C_CDNS_7230626554134 $T=423350 211195 0 0 $X=422850 $Y=210445
X170 1 VIATP_C_CDNS_7230626554134 $T=424350 211195 0 0 $X=423850 $Y=210445
X171 1 VIATP_C_CDNS_7230626554134 $T=425350 211195 0 0 $X=424850 $Y=210445
X172 1 VIATP_C_CDNS_7230626554134 $T=426350 211195 0 0 $X=425850 $Y=210445
X173 1 VIATP_C_CDNS_7230626554134 $T=427350 211195 0 0 $X=426850 $Y=210445
X174 1 VIATP_C_CDNS_7230626554134 $T=428350 211195 0 0 $X=427850 $Y=210445
X175 1 VIATP_C_CDNS_7230626554134 $T=429350 211195 0 0 $X=428850 $Y=210445
X176 1 VIATP_C_CDNS_7230626554134 $T=430350 211195 0 0 $X=429850 $Y=210445
X177 1 VIATP_C_CDNS_7230626554134 $T=431350 211195 0 0 $X=430850 $Y=210445
X178 1 VIATP_C_CDNS_7230626554134 $T=432350 211195 0 0 $X=431850 $Y=210445
X179 5 VIATP_C_CDNS_7230626554136 $T=287035 145865 0 0 $X=286535 $Y=145245
X180 5 VIATP_C_CDNS_7230626554136 $T=288035 145865 0 0 $X=287535 $Y=145245
X181 5 VIATP_C_CDNS_7230626554136 $T=289035 145865 0 0 $X=288535 $Y=145245
X182 5 VIATP_C_CDNS_7230626554136 $T=290035 145865 0 0 $X=289535 $Y=145245
X183 5 VIATP_C_CDNS_7230626554136 $T=291035 145865 0 0 $X=290535 $Y=145245
X184 5 VIATP_C_CDNS_7230626554136 $T=292035 145865 0 0 $X=291535 $Y=145245
X185 5 VIATP_C_CDNS_7230626554136 $T=293035 145865 0 0 $X=292535 $Y=145245
X186 5 VIATP_C_CDNS_7230626554136 $T=294035 145865 0 0 $X=293535 $Y=145245
X187 5 VIATP_C_CDNS_7230626554136 $T=295035 145865 0 0 $X=294535 $Y=145245
X188 5 VIATP_C_CDNS_7230626554136 $T=296035 145865 0 0 $X=295535 $Y=145245
X189 5 VIATP_C_CDNS_7230626554136 $T=395035 145865 0 0 $X=394535 $Y=145245
X190 5 VIATP_C_CDNS_7230626554136 $T=396035 145865 0 0 $X=395535 $Y=145245
X191 5 VIATP_C_CDNS_7230626554136 $T=397035 145865 0 0 $X=396535 $Y=145245
X192 5 VIATP_C_CDNS_7230626554136 $T=398035 145865 0 0 $X=397535 $Y=145245
X193 5 VIATP_C_CDNS_7230626554136 $T=399035 145865 0 0 $X=398535 $Y=145245
X194 5 VIATP_C_CDNS_7230626554136 $T=400035 145865 0 0 $X=399535 $Y=145245
X195 5 VIATP_C_CDNS_7230626554136 $T=401035 145865 0 0 $X=400535 $Y=145245
X196 5 VIATP_C_CDNS_7230626554136 $T=402035 145865 0 0 $X=401535 $Y=145245
X197 5 VIATP_C_CDNS_7230626554136 $T=403035 145865 0 0 $X=402535 $Y=145245
X198 1 VIATP_C_CDNS_7230626554136 $T=403350 182825 0 0 $X=402850 $Y=182205
X199 5 VIATP_C_CDNS_7230626554136 $T=404035 145865 0 0 $X=403535 $Y=145245
X200 1 VIATP_C_CDNS_7230626554136 $T=404350 182825 0 0 $X=403850 $Y=182205
X201 1 VIATP_C_CDNS_7230626554136 $T=406350 182825 0 0 $X=405850 $Y=182205
X202 5 VIATP_C_CDNS_7230626554136 $T=407035 145865 0 0 $X=406535 $Y=145245
X203 1 VIATP_C_CDNS_7230626554136 $T=407350 182825 0 0 $X=406850 $Y=182205
X204 5 VIATP_C_CDNS_7230626554136 $T=408035 145865 0 0 $X=407535 $Y=145245
X205 1 VIATP_C_CDNS_7230626554136 $T=408350 182825 0 0 $X=407850 $Y=182205
X206 5 VIATP_C_CDNS_7230626554136 $T=409035 145865 0 0 $X=408535 $Y=145245
X207 1 VIATP_C_CDNS_7230626554136 $T=409350 182825 0 0 $X=408850 $Y=182205
X208 5 VIATP_C_CDNS_7230626554136 $T=410035 145865 0 0 $X=409535 $Y=145245
X209 1 VIATP_C_CDNS_7230626554136 $T=410350 182825 0 0 $X=409850 $Y=182205
X210 5 VIATP_C_CDNS_7230626554136 $T=411035 145865 0 0 $X=410535 $Y=145245
X211 1 VIATP_C_CDNS_7230626554136 $T=411350 182825 0 0 $X=410850 $Y=182205
X212 5 VIATP_C_CDNS_7230626554136 $T=412035 145865 0 0 $X=411535 $Y=145245
X213 1 VIATP_C_CDNS_7230626554136 $T=412350 182825 0 0 $X=411850 $Y=182205
X214 5 VIATP_C_CDNS_7230626554136 $T=413035 145865 0 0 $X=412535 $Y=145245
X215 1 VIATP_C_CDNS_7230626554136 $T=413350 182825 0 0 $X=412850 $Y=182205
X216 5 VIATP_C_CDNS_7230626554136 $T=414035 145865 0 0 $X=413535 $Y=145245
X217 1 VIATP_C_CDNS_7230626554136 $T=414350 182825 0 0 $X=413850 $Y=182205
X218 5 VIATP_C_CDNS_7230626554136 $T=415035 117625 0 0 $X=414535 $Y=117005
X219 5 VIATP_C_CDNS_7230626554136 $T=415035 145865 0 0 $X=414535 $Y=145245
X220 1 VIATP_C_CDNS_7230626554136 $T=415350 182825 0 0 $X=414850 $Y=182205
X221 5 VIATP_C_CDNS_7230626554136 $T=416035 117625 0 0 $X=415535 $Y=117005
X222 5 VIATP_C_CDNS_7230626554136 $T=416035 145865 0 0 $X=415535 $Y=145245
X223 1 VIATP_C_CDNS_7230626554136 $T=416350 182825 0 0 $X=415850 $Y=182205
X224 5 VIATP_C_CDNS_7230626554136 $T=417035 117625 0 0 $X=416535 $Y=117005
X225 5 VIATP_C_CDNS_7230626554136 $T=417035 145865 0 0 $X=416535 $Y=145245
X226 1 VIATP_C_CDNS_7230626554136 $T=417350 182825 0 0 $X=416850 $Y=182205
X227 5 VIATP_C_CDNS_7230626554136 $T=418035 117625 0 0 $X=417535 $Y=117005
X228 5 VIATP_C_CDNS_7230626554136 $T=418035 145865 0 0 $X=417535 $Y=145245
X229 1 VIATP_C_CDNS_7230626554136 $T=418350 182825 0 0 $X=417850 $Y=182205
X230 5 VIATP_C_CDNS_7230626554136 $T=419035 117625 0 0 $X=418535 $Y=117005
X231 5 VIATP_C_CDNS_7230626554136 $T=419035 145865 0 0 $X=418535 $Y=145245
X232 1 VIATP_C_CDNS_7230626554136 $T=419350 182825 0 0 $X=418850 $Y=182205
X233 5 VIATP_C_CDNS_7230626554136 $T=420035 117625 0 0 $X=419535 $Y=117005
X234 5 VIATP_C_CDNS_7230626554136 $T=420035 145865 0 0 $X=419535 $Y=145245
X235 1 VIATP_C_CDNS_7230626554136 $T=420350 182825 0 0 $X=419850 $Y=182205
X236 5 VIATP_C_CDNS_7230626554136 $T=421035 117625 0 0 $X=420535 $Y=117005
X237 5 VIATP_C_CDNS_7230626554136 $T=421035 145865 0 0 $X=420535 $Y=145245
X238 1 VIATP_C_CDNS_7230626554136 $T=421350 182825 0 0 $X=420850 $Y=182205
X239 5 VIATP_C_CDNS_7230626554136 $T=422035 117625 0 0 $X=421535 $Y=117005
X240 5 VIATP_C_CDNS_7230626554136 $T=422035 145865 0 0 $X=421535 $Y=145245
X241 1 VIATP_C_CDNS_7230626554136 $T=422350 182825 0 0 $X=421850 $Y=182205
X242 5 VIATP_C_CDNS_7230626554136 $T=423035 117625 0 0 $X=422535 $Y=117005
X243 5 VIATP_C_CDNS_7230626554136 $T=423035 145865 0 0 $X=422535 $Y=145245
X244 1 VIATP_C_CDNS_7230626554136 $T=423350 182825 0 0 $X=422850 $Y=182205
X245 5 VIATP_C_CDNS_7230626554136 $T=424035 117625 0 0 $X=423535 $Y=117005
X246 5 VIATP_C_CDNS_7230626554136 $T=424035 145865 0 0 $X=423535 $Y=145245
X247 1 VIATP_C_CDNS_7230626554136 $T=424350 182825 0 0 $X=423850 $Y=182205
X248 5 VIATP_C_CDNS_7230626554136 $T=425035 117625 0 0 $X=424535 $Y=117005
X249 5 VIATP_C_CDNS_7230626554136 $T=425035 145865 0 0 $X=424535 $Y=145245
X250 1 VIATP_C_CDNS_7230626554136 $T=425350 182825 0 0 $X=424850 $Y=182205
X251 5 VIATP_C_CDNS_7230626554136 $T=426035 117625 0 0 $X=425535 $Y=117005
X252 5 VIATP_C_CDNS_7230626554136 $T=426035 145865 0 0 $X=425535 $Y=145245
X253 1 VIATP_C_CDNS_7230626554136 $T=426350 182825 0 0 $X=425850 $Y=182205
X254 5 VIATP_C_CDNS_7230626554136 $T=427035 117625 0 0 $X=426535 $Y=117005
X255 5 VIATP_C_CDNS_7230626554136 $T=427035 145865 0 0 $X=426535 $Y=145245
X256 1 VIATP_C_CDNS_7230626554136 $T=427350 182825 0 0 $X=426850 $Y=182205
X257 5 VIATP_C_CDNS_7230626554136 $T=428035 117625 0 0 $X=427535 $Y=117005
X258 5 VIATP_C_CDNS_7230626554136 $T=428035 145865 0 0 $X=427535 $Y=145245
X259 1 VIATP_C_CDNS_7230626554136 $T=428350 182825 0 0 $X=427850 $Y=182205
X260 5 VIATP_C_CDNS_7230626554136 $T=429035 117625 0 0 $X=428535 $Y=117005
X261 5 VIATP_C_CDNS_7230626554136 $T=429035 145865 0 0 $X=428535 $Y=145245
X262 1 VIATP_C_CDNS_7230626554136 $T=429350 182825 0 0 $X=428850 $Y=182205
X263 5 VIATP_C_CDNS_7230626554136 $T=430035 117625 0 0 $X=429535 $Y=117005
X264 5 VIATP_C_CDNS_7230626554136 $T=430035 145865 0 0 $X=429535 $Y=145245
X265 1 VIATP_C_CDNS_7230626554136 $T=430350 182825 0 0 $X=429850 $Y=182205
X266 5 VIATP_C_CDNS_7230626554136 $T=431035 117625 0 0 $X=430535 $Y=117005
X267 5 VIATP_C_CDNS_7230626554136 $T=431035 145865 0 0 $X=430535 $Y=145245
X268 1 VIATP_C_CDNS_7230626554136 $T=431350 182825 0 0 $X=430850 $Y=182205
X269 5 VIATP_C_CDNS_7230626554136 $T=432035 117625 0 0 $X=431535 $Y=117005
X270 5 VIATP_C_CDNS_7230626554136 $T=432035 145865 0 0 $X=431535 $Y=145245
X271 1 VIATP_C_CDNS_7230626554136 $T=432350 182825 0 0 $X=431850 $Y=182205
X272 5 VIATP_C_CDNS_7230626554136 $T=433035 117625 0 0 $X=432535 $Y=117005
X273 5 VIATP_C_CDNS_7230626554136 $T=433035 145865 0 0 $X=432535 $Y=145245
X274 1 VIATP_C_CDNS_7230626554137 $T=402405 182825 0 0 $X=401965 $Y=182205
X275 1 VIATP_C_CDNS_7230626554138 $T=298975 182825 0 0 $X=298100 $Y=182205
X276 1 VIATP_C_CDNS_7230626554138 $T=433725 182825 0 0 $X=432850 $Y=182205
X277 1 VIATP_C_CDNS_7230626554139 $T=298975 211195 0 0 $X=298100 $Y=210445
X278 1 VIATP_C_CDNS_7230626554139 $T=433725 211195 0 0 $X=432850 $Y=210445
X279 1 VIATP_C_CDNS_7230626554140 $T=396350 190885 0 0 $X=395850 $Y=190445
X280 1 VIATP_C_CDNS_7230626554140 $T=397350 190885 0 0 $X=396850 $Y=190445
X281 1 VIATP_C_CDNS_7230626554140 $T=398350 190885 0 0 $X=397850 $Y=190445
X282 1 VIATP_C_CDNS_7230626554140 $T=399350 190885 0 0 $X=398850 $Y=190445
X283 1 VIATP_C_CDNS_7230626554140 $T=400350 190885 0 0 $X=399850 $Y=190445
X284 1 VIATP_C_CDNS_7230626554140 $T=401350 190885 0 0 $X=400850 $Y=190445
X285 1 VIATP_C_CDNS_7230626554140 $T=402350 190885 0 0 $X=401850 $Y=190445
X286 1 VIATP_C_CDNS_7230626554142 $T=288855 191945 0 0 $X=279610 $Y=191445
X287 1 VIATP_C_CDNS_7230626554142 $T=288855 192945 0 0 $X=279610 $Y=192445
X288 1 VIATP_C_CDNS_7230626554142 $T=288855 193945 0 0 $X=279610 $Y=193445
X289 1 VIATP_C_CDNS_7230626554142 $T=288855 194945 0 0 $X=279610 $Y=194445
X290 1 VIATP_C_CDNS_7230626554142 $T=288855 195945 0 0 $X=279610 $Y=195445
X291 1 VIATP_C_CDNS_7230626554142 $T=288855 196945 0 0 $X=279610 $Y=196445
X292 1 VIATP_C_CDNS_7230626554142 $T=288855 197945 0 0 $X=279610 $Y=197445
X293 1 VIATP_C_CDNS_7230626554142 $T=288855 198945 0 0 $X=279610 $Y=198445
X294 1 VIATP_C_CDNS_7230626554142 $T=288855 199945 0 0 $X=279610 $Y=199445
X295 1 VIATP_C_CDNS_7230626554142 $T=288855 200945 0 0 $X=279610 $Y=200445
X296 1 VIATP_C_CDNS_7230626554142 $T=288855 201945 0 0 $X=279610 $Y=201445
X297 1 VIATP_C_CDNS_7230626554142 $T=288855 202945 0 0 $X=279610 $Y=202445
X298 1 VIATP_C_CDNS_7230626554142 $T=288855 203945 0 0 $X=279610 $Y=203445
X299 1 VIATP_C_CDNS_7230626554142 $T=288855 204945 0 0 $X=279610 $Y=204445
X300 5 VIATP_C_CDNS_7230626554144 $T=434275 118745 0 0 $X=433535 $Y=118245
X301 5 VIATP_C_CDNS_7230626554144 $T=434275 119745 0 0 $X=433535 $Y=119245
X302 5 VIATP_C_CDNS_7230626554144 $T=434275 120745 0 0 $X=433535 $Y=120245
X303 5 VIATP_C_CDNS_7230626554144 $T=434275 121745 0 0 $X=433535 $Y=121245
X304 5 VIATP_C_CDNS_7230626554144 $T=434275 122745 0 0 $X=433535 $Y=122245
X305 5 VIATP_C_CDNS_7230626554144 $T=434275 123745 0 0 $X=433535 $Y=123245
X306 5 VIATP_C_CDNS_7230626554144 $T=434275 124745 0 0 $X=433535 $Y=124245
X307 5 VIATP_C_CDNS_7230626554144 $T=434275 125745 0 0 $X=433535 $Y=125245
X308 5 VIATP_C_CDNS_7230626554144 $T=434275 126745 0 0 $X=433535 $Y=126245
X309 5 VIATP_C_CDNS_7230626554144 $T=434275 127745 0 0 $X=433535 $Y=127245
X310 5 VIATP_C_CDNS_7230626554144 $T=434275 128745 0 0 $X=433535 $Y=128245
X311 5 VIATP_C_CDNS_7230626554144 $T=434275 129745 0 0 $X=433535 $Y=129245
X312 5 VIATP_C_CDNS_7230626554144 $T=434275 130745 0 0 $X=433535 $Y=130245
X313 5 VIATP_C_CDNS_7230626554144 $T=434275 131745 0 0 $X=433535 $Y=131245
X314 5 VIATP_C_CDNS_7230626554144 $T=434275 132745 0 0 $X=433535 $Y=132245
X315 5 VIATP_C_CDNS_7230626554144 $T=434275 133745 0 0 $X=433535 $Y=133245
X316 5 VIATP_C_CDNS_7230626554144 $T=434275 134745 0 0 $X=433535 $Y=134245
X317 5 VIATP_C_CDNS_7230626554144 $T=434275 135745 0 0 $X=433535 $Y=135245
X318 5 VIATP_C_CDNS_7230626554144 $T=434275 136745 0 0 $X=433535 $Y=136245
X319 5 VIATP_C_CDNS_7230626554144 $T=434275 137745 0 0 $X=433535 $Y=137245
X320 5 VIATP_C_CDNS_7230626554144 $T=434275 138745 0 0 $X=433535 $Y=138245
X321 5 VIATP_C_CDNS_7230626554144 $T=434275 139745 0 0 $X=433535 $Y=139245
X322 5 VIATP_C_CDNS_7230626554144 $T=434275 140745 0 0 $X=433535 $Y=140245
X323 5 VIATP_C_CDNS_7230626554144 $T=434275 141745 0 0 $X=433535 $Y=141245
X324 5 VIATP_C_CDNS_7230626554144 $T=434275 142745 0 0 $X=433535 $Y=142245
X325 5 VIATP_C_CDNS_7230626554144 $T=434275 143745 0 0 $X=433535 $Y=143245
X326 5 VIATP_C_CDNS_7230626554144 $T=434275 144745 0 0 $X=433535 $Y=144245
X327 5 VIATP_C_CDNS_7230626554145 $T=405785 128745 0 0 $X=405515 $Y=128245
X328 5 VIATP_C_CDNS_7230626554145 $T=405785 129745 0 0 $X=405515 $Y=129245
X329 5 VIATP_C_CDNS_7230626554145 $T=405785 130745 0 0 $X=405515 $Y=130245
X330 5 VIATP_C_CDNS_7230626554145 $T=405785 131745 0 0 $X=405515 $Y=131245
X331 5 VIATP_C_CDNS_7230626554145 $T=405785 132745 0 0 $X=405515 $Y=132245
X332 5 VIATP_C_CDNS_7230626554145 $T=405785 133745 0 0 $X=405515 $Y=133245
X333 5 VIATP_C_CDNS_7230626554145 $T=405785 134745 0 0 $X=405515 $Y=134245
X334 5 VIATP_C_CDNS_7230626554145 $T=405785 135745 0 0 $X=405515 $Y=135245
X335 5 VIATP_C_CDNS_7230626554145 $T=405785 136745 0 0 $X=405515 $Y=136245
X336 5 VIATP_C_CDNS_7230626554145 $T=405785 137745 0 0 $X=405515 $Y=137245
X337 5 VIATP_C_CDNS_7230626554145 $T=405785 138745 0 0 $X=405515 $Y=138245
X338 5 VIATP_C_CDNS_7230626554145 $T=405785 139745 0 0 $X=405515 $Y=139245
X339 5 VIATP_C_CDNS_7230626554145 $T=405785 140745 0 0 $X=405515 $Y=140245
X340 5 VIATP_C_CDNS_7230626554145 $T=405785 141745 0 0 $X=405515 $Y=141245
X341 5 VIATP_C_CDNS_7230626554145 $T=405785 142745 0 0 $X=405515 $Y=142245
X342 5 VIATP_C_CDNS_7230626554145 $T=405785 143745 0 0 $X=405515 $Y=143245
X343 5 VIATP_C_CDNS_7230626554145 $T=405785 144745 0 0 $X=405515 $Y=144245
X344 5 VIATP_C_CDNS_7230626554147 $T=434275 117625 0 0 $X=433535 $Y=117005
X345 5 VIATP_C_CDNS_7230626554147 $T=434275 145865 0 0 $X=433535 $Y=145245
X346 5 VIATP_C_CDNS_7230626554149 $T=261795 145865 0 0 $X=261065 $Y=145245
X347 5 VIATP_C_CDNS_7230626554150 $T=297685 128745 0 0 $X=297415 $Y=128245
X348 5 VIATP_C_CDNS_7230626554150 $T=297685 129745 0 0 $X=297415 $Y=129245
X349 5 VIATP_C_CDNS_7230626554150 $T=297685 130745 0 0 $X=297415 $Y=130245
X350 5 VIATP_C_CDNS_7230626554150 $T=297685 131745 0 0 $X=297415 $Y=131245
X351 5 VIATP_C_CDNS_7230626554150 $T=297685 132745 0 0 $X=297415 $Y=132245
X352 5 VIATP_C_CDNS_7230626554150 $T=297685 133745 0 0 $X=297415 $Y=133245
X353 5 VIATP_C_CDNS_7230626554150 $T=297685 134745 0 0 $X=297415 $Y=134245
X354 5 VIATP_C_CDNS_7230626554150 $T=297685 135745 0 0 $X=297415 $Y=135245
X355 5 VIATP_C_CDNS_7230626554150 $T=297685 136745 0 0 $X=297415 $Y=136245
X356 5 VIATP_C_CDNS_7230626554150 $T=297685 137745 0 0 $X=297415 $Y=137245
X357 5 VIATP_C_CDNS_7230626554150 $T=297685 138745 0 0 $X=297415 $Y=138245
X358 5 VIATP_C_CDNS_7230626554150 $T=297685 139745 0 0 $X=297415 $Y=139245
X359 5 VIATP_C_CDNS_7230626554150 $T=297685 140745 0 0 $X=297415 $Y=140245
X360 5 VIATP_C_CDNS_7230626554150 $T=297685 141745 0 0 $X=297415 $Y=141245
X361 5 VIATP_C_CDNS_7230626554150 $T=297685 142745 0 0 $X=297415 $Y=142245
X362 5 VIATP_C_CDNS_7230626554150 $T=297685 143745 0 0 $X=297415 $Y=143245
X363 5 VIATP_C_CDNS_7230626554150 $T=297685 144745 0 0 $X=297415 $Y=144245
X364 5 VIATP_C_CDNS_7230626554151 $T=261795 128745 0 0 $X=261065 $Y=128245
X365 5 VIATP_C_CDNS_7230626554151 $T=261795 129745 0 0 $X=261065 $Y=129245
X366 5 VIATP_C_CDNS_7230626554151 $T=261795 130745 0 0 $X=261065 $Y=130245
X367 5 VIATP_C_CDNS_7230626554151 $T=261795 131745 0 0 $X=261065 $Y=131245
X368 5 VIATP_C_CDNS_7230626554151 $T=261795 132745 0 0 $X=261065 $Y=132245
X369 5 VIATP_C_CDNS_7230626554151 $T=261795 133745 0 0 $X=261065 $Y=133245
X370 5 VIATP_C_CDNS_7230626554151 $T=261795 134745 0 0 $X=261065 $Y=134245
X371 5 VIATP_C_CDNS_7230626554151 $T=261795 135745 0 0 $X=261065 $Y=135245
X372 5 VIATP_C_CDNS_7230626554151 $T=261795 136745 0 0 $X=261065 $Y=136245
X373 5 VIATP_C_CDNS_7230626554151 $T=261795 137745 0 0 $X=261065 $Y=137245
X374 5 VIATP_C_CDNS_7230626554151 $T=261795 138745 0 0 $X=261065 $Y=138245
X375 5 VIATP_C_CDNS_7230626554151 $T=261795 139745 0 0 $X=261065 $Y=139245
X376 5 VIATP_C_CDNS_7230626554151 $T=261795 140745 0 0 $X=261065 $Y=140245
X377 5 VIATP_C_CDNS_7230626554151 $T=261795 141745 0 0 $X=261065 $Y=141245
X378 5 VIATP_C_CDNS_7230626554151 $T=261795 142745 0 0 $X=261065 $Y=142245
X379 5 VIATP_C_CDNS_7230626554151 $T=261795 143745 0 0 $X=261065 $Y=143245
X380 5 VIATP_C_CDNS_7230626554151 $T=261795 144745 0 0 $X=261065 $Y=144245
X381 6 5 1 7 ped_CDNS_723062655411 $T=400000 176845 0 180 $X=288250 $Y=136895
X382 1 5 6 rpp1k1_3_CDNS_723062655412 $T=136055 114400 0 0 $X=132895 $Y=114180
X383 2 3 6 rpp1k1_3_CDNS_723062655416 $T=52025 148820 0 0 $X=48865 $Y=148600
X384 1 7 6 rpp1k1_3_CDNS_723062655416 $T=92050 169745 0 0 $X=88890 $Y=169525
X385 6 1 5 dpp20_CDNS_723062655418 $T=192770 173980 0 90 $X=131690 $Y=162900
X386 6 1 5 dpp20_CDNS_723062655418 $T=270135 174235 0 90 $X=209055 $Y=163155
X387 1 2 6 rpp1k1_3_CDNS_723062655419 $T=45635 170165 0 0 $X=42475 $Y=169945
X388 7 4 6 rpp1k1_3_CDNS_723062655419 $T=85700 148820 0 0 $X=82540 $Y=148600
X389 1 MASCO__X6 $T=405850 198445 0 0 $X=405850 $Y=198445
X390 1 MASCO__X6 $T=407850 198445 0 0 $X=407850 $Y=198445
X391 1 MASCO__X6 $T=409850 198445 0 0 $X=409850 $Y=198445
X392 1 MASCO__X6 $T=411850 198445 0 0 $X=411850 $Y=198445
X393 1 MASCO__X6 $T=413850 198445 0 0 $X=413850 $Y=198445
X394 5 MASCO__X6 $T=414535 133245 0 0 $X=414535 $Y=133245
X395 1 MASCO__X6 $T=415850 198445 0 0 $X=415850 $Y=198445
X396 5 MASCO__X6 $T=416535 133245 0 0 $X=416535 $Y=133245
X397 1 MASCO__X6 $T=417850 198445 0 0 $X=417850 $Y=198445
X398 5 MASCO__X6 $T=418535 133245 0 0 $X=418535 $Y=133245
X399 1 MASCO__X6 $T=419850 198445 0 0 $X=419850 $Y=198445
X400 5 MASCO__X6 $T=420535 133245 0 0 $X=420535 $Y=133245
X401 1 MASCO__X6 $T=421850 198445 0 0 $X=421850 $Y=198445
X402 5 MASCO__X6 $T=422535 133245 0 0 $X=422535 $Y=133245
X403 1 MASCO__X6 $T=423850 198445 0 0 $X=423850 $Y=198445
X404 5 MASCO__X6 $T=424535 133245 0 0 $X=424535 $Y=133245
X405 1 MASCO__X6 $T=425850 198445 0 0 $X=425850 $Y=198445
X406 5 MASCO__X6 $T=426535 133245 0 0 $X=426535 $Y=133245
X407 1 MASCO__X6 $T=427850 198445 0 0 $X=427850 $Y=198445
X408 5 MASCO__X6 $T=428535 133245 0 0 $X=428535 $Y=133245
X409 1 MASCO__X6 $T=429850 198445 0 0 $X=429850 $Y=198445
X410 5 MASCO__X6 $T=430535 133245 0 0 $X=430535 $Y=133245
X411 1 MASCO__X6 $T=431850 198445 0 0 $X=431850 $Y=198445
X412 5 MASCO__X6 $T=432535 133245 0 0 $X=432535 $Y=133245
X413 1 MASCO__X7 $T=405850 184445 0 0 $X=405850 $Y=184445
X414 1 MASCO__X7 $T=407850 184445 0 0 $X=407850 $Y=184445
X415 1 MASCO__X7 $T=409850 184445 0 0 $X=409850 $Y=184445
X416 1 MASCO__X7 $T=411850 184445 0 0 $X=411850 $Y=184445
X417 1 MASCO__X7 $T=413850 184445 0 0 $X=413850 $Y=184445
X418 5 MASCO__X7 $T=414535 119245 0 0 $X=414535 $Y=119245
X419 1 MASCO__X7 $T=415850 184445 0 0 $X=415850 $Y=184445
X420 5 MASCO__X7 $T=416535 119245 0 0 $X=416535 $Y=119245
X421 1 MASCO__X7 $T=417850 184445 0 0 $X=417850 $Y=184445
X422 5 MASCO__X7 $T=418535 119245 0 0 $X=418535 $Y=119245
X423 1 MASCO__X7 $T=419850 184445 0 0 $X=419850 $Y=184445
X424 5 MASCO__X7 $T=420535 119245 0 0 $X=420535 $Y=119245
X425 1 MASCO__X7 $T=421850 184445 0 0 $X=421850 $Y=184445
X426 5 MASCO__X7 $T=422535 119245 0 0 $X=422535 $Y=119245
X427 1 MASCO__X7 $T=423850 184445 0 0 $X=423850 $Y=184445
X428 5 MASCO__X7 $T=424535 119245 0 0 $X=424535 $Y=119245
X429 1 MASCO__X7 $T=425850 184445 0 0 $X=425850 $Y=184445
X430 5 MASCO__X7 $T=426535 119245 0 0 $X=426535 $Y=119245
X431 1 MASCO__X7 $T=427850 184445 0 0 $X=427850 $Y=184445
X432 5 MASCO__X7 $T=428535 119245 0 0 $X=428535 $Y=119245
X433 1 MASCO__X7 $T=429850 184445 0 0 $X=429850 $Y=184445
X434 5 MASCO__X7 $T=430535 119245 0 0 $X=430535 $Y=119245
X435 1 MASCO__X7 $T=431850 184445 0 0 $X=431850 $Y=184445
X436 5 MASCO__X7 $T=432535 119245 0 0 $X=432535 $Y=119245
X437 5 MASCO__X8 $T=263535 128245 0 0 $X=263535 $Y=128245
X438 5 MASCO__X8 $T=265535 128245 0 0 $X=265535 $Y=128245
X439 5 MASCO__X8 $T=267535 128245 0 0 $X=267535 $Y=128245
X440 5 MASCO__X8 $T=269535 128245 0 0 $X=269535 $Y=128245
X441 5 MASCO__X8 $T=271535 128245 0 0 $X=271535 $Y=128245
X442 5 MASCO__X8 $T=273535 128245 0 0 $X=273535 $Y=128245
X443 5 MASCO__X8 $T=275535 128245 0 0 $X=275535 $Y=128245
X444 5 MASCO__X8 $T=277535 128245 0 0 $X=277535 $Y=128245
X445 5 MASCO__X8 $T=279535 128245 0 0 $X=279535 $Y=128245
X446 5 MASCO__X8 $T=281535 128245 0 0 $X=281535 $Y=128245
X447 5 MASCO__X8 $T=283535 128245 0 0 $X=283535 $Y=128245
X448 5 MASCO__X8 $T=285535 128245 0 0 $X=285535 $Y=128245
X449 5 MASCO__X8 $T=287535 128245 0 0 $X=287535 $Y=128245
X450 5 MASCO__X8 $T=289535 128245 0 0 $X=289535 $Y=128245
X451 5 MASCO__X8 $T=291535 128245 0 0 $X=291535 $Y=128245
X452 5 MASCO__X8 $T=293535 128245 0 0 $X=293535 $Y=128245
X453 5 MASCO__X8 $T=295535 128245 0 0 $X=295535 $Y=128245
X454 5 MASCO__X8 $T=299535 128245 0 0 $X=299535 $Y=128245
X455 5 MASCO__X8 $T=301535 128245 0 0 $X=301535 $Y=128245
X456 5 MASCO__X8 $T=303535 128245 0 0 $X=303535 $Y=128245
X457 5 MASCO__X8 $T=305535 128245 0 0 $X=305535 $Y=128245
X458 5 MASCO__X8 $T=307535 128245 0 0 $X=307535 $Y=128245
X459 5 MASCO__X8 $T=309535 128245 0 0 $X=309535 $Y=128245
X460 5 MASCO__X8 $T=311535 128245 0 0 $X=311535 $Y=128245
X461 5 MASCO__X8 $T=313535 128245 0 0 $X=313535 $Y=128245
X462 5 MASCO__X8 $T=315535 128245 0 0 $X=315535 $Y=128245
X463 5 MASCO__X8 $T=317535 128245 0 0 $X=317535 $Y=128245
X464 5 MASCO__X8 $T=319535 128245 0 0 $X=319535 $Y=128245
X465 5 MASCO__X8 $T=321535 128245 0 0 $X=321535 $Y=128245
X466 5 MASCO__X8 $T=323535 128245 0 0 $X=323535 $Y=128245
X467 5 MASCO__X8 $T=325535 128245 0 0 $X=325535 $Y=128245
X468 5 MASCO__X8 $T=327535 128245 0 0 $X=327535 $Y=128245
X469 5 MASCO__X8 $T=329535 128245 0 0 $X=329535 $Y=128245
X470 5 MASCO__X8 $T=331535 128245 0 0 $X=331535 $Y=128245
X471 5 MASCO__X8 $T=333535 128245 0 0 $X=333535 $Y=128245
X472 5 MASCO__X8 $T=335535 128245 0 0 $X=335535 $Y=128245
X473 5 MASCO__X8 $T=337535 128245 0 0 $X=337535 $Y=128245
X474 5 MASCO__X8 $T=339535 128245 0 0 $X=339535 $Y=128245
X475 5 MASCO__X8 $T=341535 128245 0 0 $X=341535 $Y=128245
X476 5 MASCO__X8 $T=343535 128245 0 0 $X=343535 $Y=128245
X477 5 MASCO__X8 $T=345535 128245 0 0 $X=345535 $Y=128245
X478 5 MASCO__X8 $T=347535 128245 0 0 $X=347535 $Y=128245
X479 5 MASCO__X8 $T=349535 128245 0 0 $X=349535 $Y=128245
X480 5 MASCO__X8 $T=351535 128245 0 0 $X=351535 $Y=128245
X481 5 MASCO__X8 $T=353535 128245 0 0 $X=353535 $Y=128245
X482 5 MASCO__X8 $T=355535 128245 0 0 $X=355535 $Y=128245
X483 5 MASCO__X8 $T=357535 128245 0 0 $X=357535 $Y=128245
X484 5 MASCO__X8 $T=359535 128245 0 0 $X=359535 $Y=128245
X485 5 MASCO__X8 $T=361535 128245 0 0 $X=361535 $Y=128245
X486 5 MASCO__X8 $T=363535 128245 0 0 $X=363535 $Y=128245
X487 5 MASCO__X8 $T=365535 128245 0 0 $X=365535 $Y=128245
X488 5 MASCO__X8 $T=367535 128245 0 0 $X=367535 $Y=128245
X489 5 MASCO__X8 $T=369535 128245 0 0 $X=369535 $Y=128245
X490 5 MASCO__X8 $T=371535 128245 0 0 $X=371535 $Y=128245
X491 5 MASCO__X8 $T=373535 128245 0 0 $X=373535 $Y=128245
X492 5 MASCO__X8 $T=375535 128245 0 0 $X=375535 $Y=128245
X493 5 MASCO__X8 $T=377535 128245 0 0 $X=377535 $Y=128245
X494 5 MASCO__X8 $T=379535 128245 0 0 $X=379535 $Y=128245
X495 5 MASCO__X8 $T=381535 128245 0 0 $X=381535 $Y=128245
X496 5 MASCO__X8 $T=383535 128245 0 0 $X=383535 $Y=128245
X497 5 MASCO__X8 $T=385535 128245 0 0 $X=385535 $Y=128245
X498 5 MASCO__X8 $T=387535 128245 0 0 $X=387535 $Y=128245
X499 5 MASCO__X8 $T=389535 128245 0 0 $X=389535 $Y=128245
X500 5 MASCO__X8 $T=391535 128245 0 0 $X=391535 $Y=128245
X501 5 MASCO__X8 $T=393535 128245 0 0 $X=393535 $Y=128245
X502 5 MASCO__X8 $T=395535 128245 0 0 $X=395535 $Y=128245
X503 5 MASCO__X8 $T=397535 128245 0 0 $X=397535 $Y=128245
X504 5 MASCO__X8 $T=399535 128245 0 0 $X=399535 $Y=128245
X505 5 MASCO__X8 $T=401535 128245 0 0 $X=401535 $Y=128245
X506 1 MASCO__X8 $T=402850 183445 0 0 $X=402850 $Y=183445
X507 1 MASCO__X8 $T=402850 192445 0 0 $X=402850 $Y=192445
X508 5 MASCO__X8 $T=403535 128245 0 0 $X=403535 $Y=128245
X509 1 MASCO__X8 $T=406850 183445 0 0 $X=406850 $Y=183445
X510 1 MASCO__X8 $T=406850 192445 0 0 $X=406850 $Y=192445
X511 1 MASCO__X8 $T=406850 201445 0 0 $X=406850 $Y=201445
X512 1 MASCO__X8 $T=408850 183445 0 0 $X=408850 $Y=183445
X513 1 MASCO__X8 $T=408850 192445 0 0 $X=408850 $Y=192445
X514 1 MASCO__X8 $T=408850 201445 0 0 $X=408850 $Y=201445
X515 1 MASCO__X8 $T=410850 183445 0 0 $X=410850 $Y=183445
X516 1 MASCO__X8 $T=410850 192445 0 0 $X=410850 $Y=192445
X517 1 MASCO__X8 $T=410850 201445 0 0 $X=410850 $Y=201445
X518 1 MASCO__X8 $T=412850 183445 0 0 $X=412850 $Y=183445
X519 1 MASCO__X8 $T=412850 192445 0 0 $X=412850 $Y=192445
X520 1 MASCO__X8 $T=412850 201445 0 0 $X=412850 $Y=201445
X521 1 MASCO__X8 $T=414850 183445 0 0 $X=414850 $Y=183445
X522 1 MASCO__X8 $T=414850 192445 0 0 $X=414850 $Y=192445
X523 1 MASCO__X8 $T=414850 201445 0 0 $X=414850 $Y=201445
X524 5 MASCO__X8 $T=415535 118245 0 0 $X=415535 $Y=118245
X525 5 MASCO__X8 $T=415535 127245 0 0 $X=415535 $Y=127245
X526 5 MASCO__X8 $T=415535 136245 0 0 $X=415535 $Y=136245
X527 1 MASCO__X8 $T=416850 183445 0 0 $X=416850 $Y=183445
X528 1 MASCO__X8 $T=416850 192445 0 0 $X=416850 $Y=192445
X529 1 MASCO__X8 $T=416850 201445 0 0 $X=416850 $Y=201445
X530 5 MASCO__X8 $T=417535 118245 0 0 $X=417535 $Y=118245
X531 5 MASCO__X8 $T=417535 127245 0 0 $X=417535 $Y=127245
X532 5 MASCO__X8 $T=417535 136245 0 0 $X=417535 $Y=136245
X533 1 MASCO__X8 $T=418850 183445 0 0 $X=418850 $Y=183445
X534 1 MASCO__X8 $T=418850 192445 0 0 $X=418850 $Y=192445
X535 1 MASCO__X8 $T=418850 201445 0 0 $X=418850 $Y=201445
X536 5 MASCO__X8 $T=419535 118245 0 0 $X=419535 $Y=118245
X537 5 MASCO__X8 $T=419535 127245 0 0 $X=419535 $Y=127245
X538 5 MASCO__X8 $T=419535 136245 0 0 $X=419535 $Y=136245
X539 1 MASCO__X8 $T=420850 183445 0 0 $X=420850 $Y=183445
X540 1 MASCO__X8 $T=420850 192445 0 0 $X=420850 $Y=192445
X541 1 MASCO__X8 $T=420850 201445 0 0 $X=420850 $Y=201445
X542 5 MASCO__X8 $T=421535 118245 0 0 $X=421535 $Y=118245
X543 5 MASCO__X8 $T=421535 127245 0 0 $X=421535 $Y=127245
X544 5 MASCO__X8 $T=421535 136245 0 0 $X=421535 $Y=136245
X545 1 MASCO__X8 $T=422850 183445 0 0 $X=422850 $Y=183445
X546 1 MASCO__X8 $T=422850 192445 0 0 $X=422850 $Y=192445
X547 1 MASCO__X8 $T=422850 201445 0 0 $X=422850 $Y=201445
X548 5 MASCO__X8 $T=423535 118245 0 0 $X=423535 $Y=118245
X549 5 MASCO__X8 $T=423535 127245 0 0 $X=423535 $Y=127245
X550 5 MASCO__X8 $T=423535 136245 0 0 $X=423535 $Y=136245
X551 1 MASCO__X8 $T=424850 183445 0 0 $X=424850 $Y=183445
X552 1 MASCO__X8 $T=424850 192445 0 0 $X=424850 $Y=192445
X553 1 MASCO__X8 $T=424850 201445 0 0 $X=424850 $Y=201445
X554 5 MASCO__X8 $T=425535 118245 0 0 $X=425535 $Y=118245
X555 5 MASCO__X8 $T=425535 127245 0 0 $X=425535 $Y=127245
X556 5 MASCO__X8 $T=425535 136245 0 0 $X=425535 $Y=136245
X557 1 MASCO__X8 $T=426850 183445 0 0 $X=426850 $Y=183445
X558 1 MASCO__X8 $T=426850 192445 0 0 $X=426850 $Y=192445
X559 1 MASCO__X8 $T=426850 201445 0 0 $X=426850 $Y=201445
X560 5 MASCO__X8 $T=427535 118245 0 0 $X=427535 $Y=118245
X561 5 MASCO__X8 $T=427535 127245 0 0 $X=427535 $Y=127245
X562 5 MASCO__X8 $T=427535 136245 0 0 $X=427535 $Y=136245
X563 1 MASCO__X8 $T=428850 183445 0 0 $X=428850 $Y=183445
X564 1 MASCO__X8 $T=428850 192445 0 0 $X=428850 $Y=192445
X565 1 MASCO__X8 $T=428850 201445 0 0 $X=428850 $Y=201445
X566 5 MASCO__X8 $T=429535 118245 0 0 $X=429535 $Y=118245
X567 5 MASCO__X8 $T=429535 127245 0 0 $X=429535 $Y=127245
X568 5 MASCO__X8 $T=429535 136245 0 0 $X=429535 $Y=136245
X569 1 MASCO__X8 $T=430850 183445 0 0 $X=430850 $Y=183445
X570 1 MASCO__X8 $T=430850 192445 0 0 $X=430850 $Y=192445
X571 1 MASCO__X8 $T=430850 201445 0 0 $X=430850 $Y=201445
X572 5 MASCO__X8 $T=431535 118245 0 0 $X=431535 $Y=118245
X573 5 MASCO__X8 $T=431535 127245 0 0 $X=431535 $Y=127245
X574 5 MASCO__X8 $T=431535 136245 0 0 $X=431535 $Y=136245
X575 5 MASCO__X9 $T=263535 137245 0 0 $X=263535 $Y=137245
X576 5 MASCO__X9 $T=265535 137245 0 0 $X=265535 $Y=137245
X577 5 MASCO__X9 $T=267535 137245 0 0 $X=267535 $Y=137245
X578 5 MASCO__X9 $T=269535 137245 0 0 $X=269535 $Y=137245
X579 5 MASCO__X9 $T=271535 137245 0 0 $X=271535 $Y=137245
X580 5 MASCO__X9 $T=273535 137245 0 0 $X=273535 $Y=137245
X581 5 MASCO__X9 $T=275535 137245 0 0 $X=275535 $Y=137245
X582 5 MASCO__X9 $T=277535 137245 0 0 $X=277535 $Y=137245
X583 5 MASCO__X9 $T=279535 137245 0 0 $X=279535 $Y=137245
X584 5 MASCO__X9 $T=281535 137245 0 0 $X=281535 $Y=137245
X585 5 MASCO__X9 $T=283535 137245 0 0 $X=283535 $Y=137245
X586 5 MASCO__X9 $T=285535 137245 0 0 $X=285535 $Y=137245
X587 5 MASCO__X9 $T=287535 137245 0 0 $X=287535 $Y=137245
X588 5 MASCO__X9 $T=289535 137245 0 0 $X=289535 $Y=137245
X589 5 MASCO__X9 $T=291535 137245 0 0 $X=291535 $Y=137245
X590 5 MASCO__X9 $T=293535 137245 0 0 $X=293535 $Y=137245
X591 5 MASCO__X9 $T=295535 137245 0 0 $X=295535 $Y=137245
X592 5 MASCO__X9 $T=299535 137245 0 0 $X=299535 $Y=137245
X593 5 MASCO__X9 $T=301535 137245 0 0 $X=301535 $Y=137245
X594 5 MASCO__X9 $T=303535 137245 0 0 $X=303535 $Y=137245
X595 5 MASCO__X9 $T=305535 137245 0 0 $X=305535 $Y=137245
X596 5 MASCO__X9 $T=307535 137245 0 0 $X=307535 $Y=137245
X597 5 MASCO__X9 $T=309535 137245 0 0 $X=309535 $Y=137245
X598 5 MASCO__X9 $T=311535 137245 0 0 $X=311535 $Y=137245
X599 5 MASCO__X9 $T=313535 137245 0 0 $X=313535 $Y=137245
X600 5 MASCO__X9 $T=315535 137245 0 0 $X=315535 $Y=137245
X601 5 MASCO__X9 $T=317535 137245 0 0 $X=317535 $Y=137245
X602 5 MASCO__X9 $T=319535 137245 0 0 $X=319535 $Y=137245
X603 5 MASCO__X9 $T=321535 137245 0 0 $X=321535 $Y=137245
X604 5 MASCO__X9 $T=323535 137245 0 0 $X=323535 $Y=137245
X605 5 MASCO__X9 $T=325535 137245 0 0 $X=325535 $Y=137245
X606 5 MASCO__X9 $T=327535 137245 0 0 $X=327535 $Y=137245
X607 5 MASCO__X9 $T=329535 137245 0 0 $X=329535 $Y=137245
X608 5 MASCO__X9 $T=331535 137245 0 0 $X=331535 $Y=137245
X609 5 MASCO__X9 $T=333535 137245 0 0 $X=333535 $Y=137245
X610 5 MASCO__X9 $T=335535 137245 0 0 $X=335535 $Y=137245
X611 5 MASCO__X9 $T=337535 137245 0 0 $X=337535 $Y=137245
X612 5 MASCO__X9 $T=339535 137245 0 0 $X=339535 $Y=137245
X613 5 MASCO__X9 $T=341535 137245 0 0 $X=341535 $Y=137245
X614 5 MASCO__X9 $T=343535 137245 0 0 $X=343535 $Y=137245
X615 5 MASCO__X9 $T=345535 137245 0 0 $X=345535 $Y=137245
X616 5 MASCO__X9 $T=347535 137245 0 0 $X=347535 $Y=137245
X617 5 MASCO__X9 $T=349535 137245 0 0 $X=349535 $Y=137245
X618 5 MASCO__X9 $T=351535 137245 0 0 $X=351535 $Y=137245
X619 5 MASCO__X9 $T=353535 137245 0 0 $X=353535 $Y=137245
X620 5 MASCO__X9 $T=355535 137245 0 0 $X=355535 $Y=137245
X621 5 MASCO__X9 $T=357535 137245 0 0 $X=357535 $Y=137245
X622 5 MASCO__X9 $T=359535 137245 0 0 $X=359535 $Y=137245
X623 5 MASCO__X9 $T=361535 137245 0 0 $X=361535 $Y=137245
X624 5 MASCO__X9 $T=363535 137245 0 0 $X=363535 $Y=137245
X625 5 MASCO__X9 $T=365535 137245 0 0 $X=365535 $Y=137245
X626 5 MASCO__X9 $T=367535 137245 0 0 $X=367535 $Y=137245
X627 5 MASCO__X9 $T=369535 137245 0 0 $X=369535 $Y=137245
X628 5 MASCO__X9 $T=371535 137245 0 0 $X=371535 $Y=137245
X629 5 MASCO__X9 $T=373535 137245 0 0 $X=373535 $Y=137245
X630 5 MASCO__X9 $T=375535 137245 0 0 $X=375535 $Y=137245
X631 5 MASCO__X9 $T=377535 137245 0 0 $X=377535 $Y=137245
X632 5 MASCO__X9 $T=379535 137245 0 0 $X=379535 $Y=137245
X633 5 MASCO__X9 $T=381535 137245 0 0 $X=381535 $Y=137245
X634 5 MASCO__X9 $T=383535 137245 0 0 $X=383535 $Y=137245
X635 5 MASCO__X9 $T=385535 137245 0 0 $X=385535 $Y=137245
X636 5 MASCO__X9 $T=387535 137245 0 0 $X=387535 $Y=137245
X637 5 MASCO__X9 $T=389535 137245 0 0 $X=389535 $Y=137245
X638 5 MASCO__X9 $T=391535 137245 0 0 $X=391535 $Y=137245
X639 5 MASCO__X9 $T=393535 137245 0 0 $X=393535 $Y=137245
X640 5 MASCO__X9 $T=395535 137245 0 0 $X=395535 $Y=137245
X641 5 MASCO__X9 $T=397535 137245 0 0 $X=397535 $Y=137245
X642 5 MASCO__X9 $T=399535 137245 0 0 $X=399535 $Y=137245
X643 5 MASCO__X9 $T=401535 137245 0 0 $X=401535 $Y=137245
X644 5 MASCO__X9 $T=403535 137245 0 0 $X=403535 $Y=137245
X645 5 MASCO__X9 $T=407535 137245 0 0 $X=407535 $Y=137245
X646 5 MASCO__X9 $T=409535 137245 0 0 $X=409535 $Y=137245
X647 5 MASCO__X9 $T=411535 137245 0 0 $X=411535 $Y=137245
X648 5 MASCO__X9 $T=413535 137245 0 0 $X=413535 $Y=137245
X649 5 MASCO__X10 $T=262535 129245 0 0 $X=262535 $Y=129245
X650 5 MASCO__X10 $T=264535 129245 0 0 $X=264535 $Y=129245
X651 5 MASCO__X10 $T=266535 129245 0 0 $X=266535 $Y=129245
X652 5 MASCO__X10 $T=268535 129245 0 0 $X=268535 $Y=129245
X653 5 MASCO__X10 $T=270535 129245 0 0 $X=270535 $Y=129245
X654 5 MASCO__X10 $T=272535 129245 0 0 $X=272535 $Y=129245
X655 5 MASCO__X10 $T=274535 129245 0 0 $X=274535 $Y=129245
X656 5 MASCO__X10 $T=276535 129245 0 0 $X=276535 $Y=129245
X657 5 MASCO__X10 $T=278535 129245 0 0 $X=278535 $Y=129245
X658 5 MASCO__X10 $T=280535 129245 0 0 $X=280535 $Y=129245
X659 5 MASCO__X10 $T=282535 129245 0 0 $X=282535 $Y=129245
X660 5 MASCO__X10 $T=284535 129245 0 0 $X=284535 $Y=129245
X661 5 MASCO__X10 $T=286535 129245 0 0 $X=286535 $Y=129245
X662 5 MASCO__X10 $T=288535 129245 0 0 $X=288535 $Y=129245
X663 5 MASCO__X10 $T=290535 129245 0 0 $X=290535 $Y=129245
X664 5 MASCO__X10 $T=292535 129245 0 0 $X=292535 $Y=129245
X665 5 MASCO__X10 $T=294535 129245 0 0 $X=294535 $Y=129245
X666 5 MASCO__X10 $T=298535 129245 0 0 $X=298535 $Y=129245
X667 5 MASCO__X10 $T=300535 129245 0 0 $X=300535 $Y=129245
X668 5 MASCO__X10 $T=302535 129245 0 0 $X=302535 $Y=129245
X669 5 MASCO__X10 $T=304535 129245 0 0 $X=304535 $Y=129245
X670 5 MASCO__X10 $T=306535 129245 0 0 $X=306535 $Y=129245
X671 5 MASCO__X10 $T=308535 129245 0 0 $X=308535 $Y=129245
X672 5 MASCO__X10 $T=310535 129245 0 0 $X=310535 $Y=129245
X673 5 MASCO__X10 $T=312535 129245 0 0 $X=312535 $Y=129245
X674 5 MASCO__X10 $T=314535 129245 0 0 $X=314535 $Y=129245
X675 5 MASCO__X10 $T=316535 129245 0 0 $X=316535 $Y=129245
X676 5 MASCO__X10 $T=318535 129245 0 0 $X=318535 $Y=129245
X677 5 MASCO__X10 $T=320535 129245 0 0 $X=320535 $Y=129245
X678 5 MASCO__X10 $T=322535 129245 0 0 $X=322535 $Y=129245
X679 5 MASCO__X10 $T=324535 129245 0 0 $X=324535 $Y=129245
X680 5 MASCO__X10 $T=326535 129245 0 0 $X=326535 $Y=129245
X681 5 MASCO__X10 $T=328535 129245 0 0 $X=328535 $Y=129245
X682 5 MASCO__X10 $T=330535 129245 0 0 $X=330535 $Y=129245
X683 5 MASCO__X10 $T=332535 129245 0 0 $X=332535 $Y=129245
X684 5 MASCO__X10 $T=334535 129245 0 0 $X=334535 $Y=129245
X685 5 MASCO__X10 $T=336535 129245 0 0 $X=336535 $Y=129245
X686 5 MASCO__X10 $T=338535 129245 0 0 $X=338535 $Y=129245
X687 5 MASCO__X10 $T=340535 129245 0 0 $X=340535 $Y=129245
X688 5 MASCO__X10 $T=342535 129245 0 0 $X=342535 $Y=129245
X689 5 MASCO__X10 $T=344535 129245 0 0 $X=344535 $Y=129245
X690 5 MASCO__X10 $T=346535 129245 0 0 $X=346535 $Y=129245
X691 5 MASCO__X10 $T=348535 129245 0 0 $X=348535 $Y=129245
X692 5 MASCO__X10 $T=350535 129245 0 0 $X=350535 $Y=129245
X693 5 MASCO__X10 $T=352535 129245 0 0 $X=352535 $Y=129245
X694 5 MASCO__X10 $T=354535 129245 0 0 $X=354535 $Y=129245
X695 5 MASCO__X10 $T=356535 129245 0 0 $X=356535 $Y=129245
X696 5 MASCO__X10 $T=358535 129245 0 0 $X=358535 $Y=129245
X697 5 MASCO__X10 $T=360535 129245 0 0 $X=360535 $Y=129245
X698 5 MASCO__X10 $T=362535 129245 0 0 $X=362535 $Y=129245
X699 5 MASCO__X10 $T=364535 129245 0 0 $X=364535 $Y=129245
X700 5 MASCO__X10 $T=366535 129245 0 0 $X=366535 $Y=129245
X701 5 MASCO__X10 $T=368535 129245 0 0 $X=368535 $Y=129245
X702 5 MASCO__X10 $T=370535 129245 0 0 $X=370535 $Y=129245
X703 5 MASCO__X10 $T=372535 129245 0 0 $X=372535 $Y=129245
X704 5 MASCO__X10 $T=374535 129245 0 0 $X=374535 $Y=129245
X705 5 MASCO__X10 $T=376535 129245 0 0 $X=376535 $Y=129245
X706 5 MASCO__X10 $T=378535 129245 0 0 $X=378535 $Y=129245
X707 5 MASCO__X10 $T=380535 129245 0 0 $X=380535 $Y=129245
X708 5 MASCO__X10 $T=382535 129245 0 0 $X=382535 $Y=129245
X709 5 MASCO__X10 $T=384535 129245 0 0 $X=384535 $Y=129245
X710 5 MASCO__X10 $T=386535 129245 0 0 $X=386535 $Y=129245
X711 5 MASCO__X10 $T=388535 129245 0 0 $X=388535 $Y=129245
X712 5 MASCO__X10 $T=390535 129245 0 0 $X=390535 $Y=129245
X713 5 MASCO__X10 $T=392535 129245 0 0 $X=392535 $Y=129245
X714 5 MASCO__X10 $T=394535 129245 0 0 $X=394535 $Y=129245
X715 5 MASCO__X10 $T=396535 129245 0 0 $X=396535 $Y=129245
X716 5 MASCO__X10 $T=398535 129245 0 0 $X=398535 $Y=129245
X717 5 MASCO__X10 $T=400535 129245 0 0 $X=400535 $Y=129245
X718 5 MASCO__X10 $T=402535 129245 0 0 $X=402535 $Y=129245
X719 5 MASCO__X10 $T=406535 129245 0 0 $X=406535 $Y=129245
X720 5 MASCO__X10 $T=408535 129245 0 0 $X=408535 $Y=129245
X721 5 MASCO__X10 $T=410535 129245 0 0 $X=410535 $Y=129245
X722 5 MASCO__X10 $T=412535 129245 0 0 $X=412535 $Y=129245
X723 1 MASCO__X12 $T=300850 191445 0 0 $X=300850 $Y=191445
X724 1 MASCO__X12 $T=302850 191445 0 0 $X=302850 $Y=191445
X725 1 MASCO__X12 $T=304850 191445 0 0 $X=304850 $Y=191445
X726 1 MASCO__X12 $T=306850 191445 0 0 $X=306850 $Y=191445
X727 1 MASCO__X12 $T=308850 191445 0 0 $X=308850 $Y=191445
X728 1 MASCO__X12 $T=310850 191445 0 0 $X=310850 $Y=191445
X729 1 MASCO__X12 $T=312850 191445 0 0 $X=312850 $Y=191445
X730 1 MASCO__X12 $T=314850 191445 0 0 $X=314850 $Y=191445
X731 1 MASCO__X12 $T=316850 191445 0 0 $X=316850 $Y=191445
X732 1 MASCO__X12 $T=318850 191445 0 0 $X=318850 $Y=191445
X733 1 MASCO__X12 $T=320850 191445 0 0 $X=320850 $Y=191445
X734 1 MASCO__X12 $T=322850 191445 0 0 $X=322850 $Y=191445
X735 1 MASCO__X12 $T=324850 191445 0 0 $X=324850 $Y=191445
X736 1 MASCO__X12 $T=326850 191445 0 0 $X=326850 $Y=191445
X737 1 MASCO__X12 $T=328850 191445 0 0 $X=328850 $Y=191445
X738 1 MASCO__X12 $T=330850 191445 0 0 $X=330850 $Y=191445
X739 1 MASCO__X12 $T=332850 191445 0 0 $X=332850 $Y=191445
X740 1 MASCO__X12 $T=334850 191445 0 0 $X=334850 $Y=191445
X741 1 MASCO__X12 $T=336850 191445 0 0 $X=336850 $Y=191445
X742 1 MASCO__X12 $T=338850 191445 0 0 $X=338850 $Y=191445
X743 1 MASCO__X12 $T=340850 191445 0 0 $X=340850 $Y=191445
X744 1 MASCO__X12 $T=342850 191445 0 0 $X=342850 $Y=191445
X745 1 MASCO__X12 $T=344850 191445 0 0 $X=344850 $Y=191445
X746 1 MASCO__X12 $T=346850 191445 0 0 $X=346850 $Y=191445
X747 1 MASCO__X12 $T=348850 191445 0 0 $X=348850 $Y=191445
X748 1 MASCO__X12 $T=350850 191445 0 0 $X=350850 $Y=191445
X749 1 MASCO__X12 $T=352850 191445 0 0 $X=352850 $Y=191445
X750 1 MASCO__X12 $T=354850 191445 0 0 $X=354850 $Y=191445
X751 1 MASCO__X12 $T=356850 191445 0 0 $X=356850 $Y=191445
X752 1 MASCO__X12 $T=358850 191445 0 0 $X=358850 $Y=191445
X753 1 MASCO__X12 $T=360850 191445 0 0 $X=360850 $Y=191445
X754 1 MASCO__X12 $T=362850 191445 0 0 $X=362850 $Y=191445
X755 1 MASCO__X12 $T=364850 191445 0 0 $X=364850 $Y=191445
X756 1 MASCO__X12 $T=366850 191445 0 0 $X=366850 $Y=191445
X757 1 MASCO__X12 $T=368850 191445 0 0 $X=368850 $Y=191445
X758 1 MASCO__X12 $T=370850 191445 0 0 $X=370850 $Y=191445
X759 1 MASCO__X12 $T=372850 191445 0 0 $X=372850 $Y=191445
X760 1 MASCO__X12 $T=374850 191445 0 0 $X=374850 $Y=191445
X761 1 MASCO__X12 $T=376850 191445 0 0 $X=376850 $Y=191445
X762 1 MASCO__X12 $T=378850 191445 0 0 $X=378850 $Y=191445
X763 1 MASCO__X12 $T=380850 191445 0 0 $X=380850 $Y=191445
X764 1 MASCO__X12 $T=382850 191445 0 0 $X=382850 $Y=191445
X765 1 MASCO__X12 $T=384850 191445 0 0 $X=384850 $Y=191445
X766 1 MASCO__X12 $T=386850 191445 0 0 $X=386850 $Y=191445
X767 1 MASCO__X12 $T=388850 191445 0 0 $X=388850 $Y=191445
X768 1 MASCO__X12 $T=390850 191445 0 0 $X=390850 $Y=191445
X769 1 MASCO__X12 $T=392850 191445 0 0 $X=392850 $Y=191445
X770 1 MASCO__X12 $T=394850 191445 0 0 $X=394850 $Y=191445
X771 1 MASCO__X12 $T=396850 191445 0 0 $X=396850 $Y=191445
X772 1 MASCO__X12 $T=398850 191445 0 0 $X=398850 $Y=191445
X773 1 MASCO__X12 $T=400850 191445 0 0 $X=400850 $Y=191445
X774 1 MASCO__X13 $T=300850 183445 0 0 $X=300850 $Y=183445
X775 1 MASCO__X13 $T=302850 183445 0 0 $X=302850 $Y=183445
X776 1 MASCO__X13 $T=304850 183445 0 0 $X=304850 $Y=183445
X777 1 MASCO__X13 $T=306850 183445 0 0 $X=306850 $Y=183445
X778 1 MASCO__X13 $T=308850 183445 0 0 $X=308850 $Y=183445
X779 1 MASCO__X13 $T=310850 183445 0 0 $X=310850 $Y=183445
X780 1 MASCO__X13 $T=312850 183445 0 0 $X=312850 $Y=183445
X781 1 MASCO__X13 $T=314850 183445 0 0 $X=314850 $Y=183445
X782 1 MASCO__X13 $T=316850 183445 0 0 $X=316850 $Y=183445
X783 1 MASCO__X13 $T=318850 183445 0 0 $X=318850 $Y=183445
X784 1 MASCO__X13 $T=320850 183445 0 0 $X=320850 $Y=183445
X785 1 MASCO__X13 $T=322850 183445 0 0 $X=322850 $Y=183445
X786 1 MASCO__X13 $T=324850 183445 0 0 $X=324850 $Y=183445
X787 1 MASCO__X13 $T=326850 183445 0 0 $X=326850 $Y=183445
X788 1 MASCO__X13 $T=328850 183445 0 0 $X=328850 $Y=183445
X789 1 MASCO__X13 $T=330850 183445 0 0 $X=330850 $Y=183445
X790 1 MASCO__X13 $T=332850 183445 0 0 $X=332850 $Y=183445
X791 1 MASCO__X13 $T=334850 183445 0 0 $X=334850 $Y=183445
X792 1 MASCO__X13 $T=336850 183445 0 0 $X=336850 $Y=183445
X793 1 MASCO__X13 $T=338850 183445 0 0 $X=338850 $Y=183445
X794 1 MASCO__X13 $T=340850 183445 0 0 $X=340850 $Y=183445
X795 1 MASCO__X13 $T=342850 183445 0 0 $X=342850 $Y=183445
X796 1 MASCO__X13 $T=344850 183445 0 0 $X=344850 $Y=183445
X797 1 MASCO__X13 $T=346850 183445 0 0 $X=346850 $Y=183445
X798 1 MASCO__X13 $T=348850 183445 0 0 $X=348850 $Y=183445
X799 1 MASCO__X13 $T=350850 183445 0 0 $X=350850 $Y=183445
X800 1 MASCO__X13 $T=352850 183445 0 0 $X=352850 $Y=183445
X801 1 MASCO__X13 $T=354850 183445 0 0 $X=354850 $Y=183445
X802 1 MASCO__X13 $T=356850 183445 0 0 $X=356850 $Y=183445
X803 1 MASCO__X13 $T=358850 183445 0 0 $X=358850 $Y=183445
X804 1 MASCO__X13 $T=360850 183445 0 0 $X=360850 $Y=183445
X805 1 MASCO__X13 $T=362850 183445 0 0 $X=362850 $Y=183445
X806 1 MASCO__X13 $T=364850 183445 0 0 $X=364850 $Y=183445
X807 1 MASCO__X13 $T=366850 183445 0 0 $X=366850 $Y=183445
X808 1 MASCO__X13 $T=368850 183445 0 0 $X=368850 $Y=183445
X809 1 MASCO__X13 $T=370850 183445 0 0 $X=370850 $Y=183445
X810 1 MASCO__X13 $T=372850 183445 0 0 $X=372850 $Y=183445
X811 1 MASCO__X13 $T=374850 183445 0 0 $X=374850 $Y=183445
X812 1 MASCO__X13 $T=376850 183445 0 0 $X=376850 $Y=183445
X813 1 MASCO__X13 $T=378850 183445 0 0 $X=378850 $Y=183445
X814 1 MASCO__X13 $T=380850 183445 0 0 $X=380850 $Y=183445
X815 1 MASCO__X13 $T=382850 183445 0 0 $X=382850 $Y=183445
X816 1 MASCO__X13 $T=384850 183445 0 0 $X=384850 $Y=183445
X817 1 MASCO__X13 $T=386850 183445 0 0 $X=386850 $Y=183445
X818 1 MASCO__X13 $T=388850 183445 0 0 $X=388850 $Y=183445
X819 1 MASCO__X13 $T=390850 183445 0 0 $X=390850 $Y=183445
X820 1 MASCO__X13 $T=392850 183445 0 0 $X=392850 $Y=183445
X821 1 MASCO__X13 $T=394850 183445 0 0 $X=394850 $Y=183445
X822 1 MASCO__X13 $T=396850 183445 0 0 $X=396850 $Y=183445
X823 1 MASCO__X13 $T=398850 183445 0 0 $X=398850 $Y=183445
X824 1 MASCO__X13 $T=400850 183445 0 0 $X=400850 $Y=183445
X825 1 MASCO__Y15 $T=299850 190445 0 0 $X=299850 $Y=190445
X826 1 MASCO__Y15 $T=311850 190445 0 0 $X=311850 $Y=190445
X827 1 MASCO__Y15 $T=323850 190445 0 0 $X=323850 $Y=190445
X828 1 MASCO__Y15 $T=335850 190445 0 0 $X=335850 $Y=190445
X829 1 MASCO__Y15 $T=347850 190445 0 0 $X=347850 $Y=190445
X830 1 MASCO__Y15 $T=359850 190445 0 0 $X=359850 $Y=190445
X831 1 MASCO__Y15 $T=371850 190445 0 0 $X=371850 $Y=190445
X832 1 MASCO__Y15 $T=383850 190445 0 0 $X=383850 $Y=190445
X833 1 MASCO__Y16 $T=299850 192445 0 0 $X=299850 $Y=192445
X834 1 MASCO__Y16 $T=307850 192445 0 0 $X=307850 $Y=192445
X835 1 MASCO__Y16 $T=315850 192445 0 0 $X=315850 $Y=192445
X836 1 MASCO__Y16 $T=323850 192445 0 0 $X=323850 $Y=192445
X837 1 MASCO__Y16 $T=331850 192445 0 0 $X=331850 $Y=192445
X838 1 MASCO__Y16 $T=339850 192445 0 0 $X=339850 $Y=192445
X839 1 MASCO__Y16 $T=347850 192445 0 0 $X=347850 $Y=192445
X840 1 MASCO__Y16 $T=355850 192445 0 0 $X=355850 $Y=192445
X841 1 MASCO__Y16 $T=363850 192445 0 0 $X=363850 $Y=192445
X842 1 MASCO__Y16 $T=371850 192445 0 0 $X=371850 $Y=192445
X843 1 MASCO__Y16 $T=379850 192445 0 0 $X=379850 $Y=192445
X844 1 MASCO__Y16 $T=387850 192445 0 0 $X=387850 $Y=192445
X845 1 MASCO__Y16 $T=395850 192445 0 0 $X=395850 $Y=192445
X846 1 MASCO__Y17 $T=299850 182205 0 0 $X=299850 $Y=182205
X847 1 MASCO__Y17 $T=305850 182205 0 0 $X=305850 $Y=182205
X848 1 MASCO__Y17 $T=311850 182205 0 0 $X=311850 $Y=182205
X849 1 MASCO__Y17 $T=317850 182205 0 0 $X=317850 $Y=182205
X850 1 MASCO__Y17 $T=323850 182205 0 0 $X=323850 $Y=182205
X851 1 MASCO__Y17 $T=329850 182205 0 0 $X=329850 $Y=182205
X852 1 MASCO__Y17 $T=335850 182205 0 0 $X=335850 $Y=182205
X853 1 MASCO__Y17 $T=341850 182205 0 0 $X=341850 $Y=182205
X854 1 MASCO__Y17 $T=347850 182205 0 0 $X=347850 $Y=182205
X855 1 MASCO__Y17 $T=353850 182205 0 0 $X=353850 $Y=182205
X856 1 MASCO__Y17 $T=359850 182205 0 0 $X=359850 $Y=182205
X857 1 MASCO__Y17 $T=365850 182205 0 0 $X=365850 $Y=182205
X858 1 MASCO__Y17 $T=371850 182205 0 0 $X=371850 $Y=182205
X859 1 MASCO__Y17 $T=377850 182205 0 0 $X=377850 $Y=182205
X860 1 MASCO__Y17 $T=383850 182205 0 0 $X=383850 $Y=182205
X861 1 MASCO__Y17 $T=389850 182205 0 0 $X=389850 $Y=182205
X862 1 MASCO__Y17 $T=395850 182205 0 0 $X=395850 $Y=182205
X863 5 MASCO__Y18 $T=262535 145245 0 0 $X=262535 $Y=145245
X864 5 MASCO__Y18 $T=274535 145245 0 0 $X=274535 $Y=145245
X865 5 MASCO__Y18 $T=298535 145245 0 0 $X=298535 $Y=145245
X866 5 MASCO__Y18 $T=310535 145245 0 0 $X=310535 $Y=145245
X867 5 MASCO__Y18 $T=322535 145245 0 0 $X=322535 $Y=145245
X868 5 MASCO__Y18 $T=334535 145245 0 0 $X=334535 $Y=145245
X869 5 MASCO__Y18 $T=346535 145245 0 0 $X=346535 $Y=145245
X870 5 MASCO__Y18 $T=358535 145245 0 0 $X=358535 $Y=145245
X871 5 MASCO__Y18 $T=370535 145245 0 0 $X=370535 $Y=145245
X872 5 MASCO__Y18 $T=382535 145245 0 0 $X=382535 $Y=145245
X873 1 MASCO__Y19 $T=300850 201445 0 0 $X=300850 $Y=201445
X874 1 MASCO__Y19 $T=308850 201445 0 0 $X=308850 $Y=201445
X875 1 MASCO__Y19 $T=316850 201445 0 0 $X=316850 $Y=201445
X876 1 MASCO__Y19 $T=324850 201445 0 0 $X=324850 $Y=201445
X877 1 MASCO__Y19 $T=332850 201445 0 0 $X=332850 $Y=201445
X878 1 MASCO__Y19 $T=340850 201445 0 0 $X=340850 $Y=201445
X879 1 MASCO__Y19 $T=348850 201445 0 0 $X=348850 $Y=201445
X880 1 MASCO__Y19 $T=356850 201445 0 0 $X=356850 $Y=201445
X881 1 MASCO__Y19 $T=364850 201445 0 0 $X=364850 $Y=201445
X882 1 MASCO__Y19 $T=372850 201445 0 0 $X=372850 $Y=201445
X883 1 MASCO__Y19 $T=380850 201445 0 0 $X=380850 $Y=201445
X884 1 MASCO__Y19 $T=388850 201445 0 0 $X=388850 $Y=201445
X885 1 MASCO__Y19 $T=396850 201445 0 0 $X=396850 $Y=201445
X886 5 MASCO__Y19 $T=407535 128245 0 0 $X=407535 $Y=128245
X887 1 MASCO__Y20 $T=299850 210445 0 0 $X=299850 $Y=210445
X888 1 MASCO__Y20 $T=307850 210445 0 0 $X=307850 $Y=210445
X889 1 MASCO__Y20 $T=315850 210445 0 0 $X=315850 $Y=210445
X890 1 MASCO__Y20 $T=323850 210445 0 0 $X=323850 $Y=210445
X891 1 MASCO__Y20 $T=331850 210445 0 0 $X=331850 $Y=210445
X892 1 MASCO__Y20 $T=339850 210445 0 0 $X=339850 $Y=210445
X893 1 MASCO__Y20 $T=347850 210445 0 0 $X=347850 $Y=210445
X894 1 MASCO__Y20 $T=355850 210445 0 0 $X=355850 $Y=210445
X895 1 MASCO__Y20 $T=363850 210445 0 0 $X=363850 $Y=210445
X896 1 MASCO__Y20 $T=371850 210445 0 0 $X=371850 $Y=210445
X897 1 MASCO__Y20 $T=379850 210445 0 0 $X=379850 $Y=210445
X898 1 MASCO__Y20 $T=387850 210445 0 0 $X=387850 $Y=210445
X899 1 MASCO__Y20 $T=395850 210445 0 0 $X=395850 $Y=210445
X900 1 MASCO__Y21 $T=299850 184445 0 0 $X=299850 $Y=184445
X901 1 MASCO__Y21 $T=299850 186445 0 0 $X=299850 $Y=186445
X902 1 MASCO__Y21 $T=299850 188445 0 0 $X=299850 $Y=188445
X903 1 MASCO__Y21 $T=307850 184445 0 0 $X=307850 $Y=184445
X904 1 MASCO__Y21 $T=307850 186445 0 0 $X=307850 $Y=186445
X905 1 MASCO__Y21 $T=307850 188445 0 0 $X=307850 $Y=188445
X906 1 MASCO__Y21 $T=315850 184445 0 0 $X=315850 $Y=184445
X907 1 MASCO__Y21 $T=315850 186445 0 0 $X=315850 $Y=186445
X908 1 MASCO__Y21 $T=315850 188445 0 0 $X=315850 $Y=188445
X909 1 MASCO__Y21 $T=323850 184445 0 0 $X=323850 $Y=184445
X910 1 MASCO__Y21 $T=323850 186445 0 0 $X=323850 $Y=186445
X911 1 MASCO__Y21 $T=323850 188445 0 0 $X=323850 $Y=188445
X912 1 MASCO__Y21 $T=331850 184445 0 0 $X=331850 $Y=184445
X913 1 MASCO__Y21 $T=331850 186445 0 0 $X=331850 $Y=186445
X914 1 MASCO__Y21 $T=331850 188445 0 0 $X=331850 $Y=188445
X915 1 MASCO__Y21 $T=339850 184445 0 0 $X=339850 $Y=184445
X916 1 MASCO__Y21 $T=339850 186445 0 0 $X=339850 $Y=186445
X917 1 MASCO__Y21 $T=339850 188445 0 0 $X=339850 $Y=188445
X918 1 MASCO__Y21 $T=347850 184445 0 0 $X=347850 $Y=184445
X919 1 MASCO__Y21 $T=347850 186445 0 0 $X=347850 $Y=186445
X920 1 MASCO__Y21 $T=347850 188445 0 0 $X=347850 $Y=188445
X921 1 MASCO__Y21 $T=355850 184445 0 0 $X=355850 $Y=184445
X922 1 MASCO__Y21 $T=355850 186445 0 0 $X=355850 $Y=186445
X923 1 MASCO__Y21 $T=355850 188445 0 0 $X=355850 $Y=188445
X924 1 MASCO__Y21 $T=363850 184445 0 0 $X=363850 $Y=184445
X925 1 MASCO__Y21 $T=363850 186445 0 0 $X=363850 $Y=186445
X926 1 MASCO__Y21 $T=363850 188445 0 0 $X=363850 $Y=188445
X927 1 MASCO__Y21 $T=371850 184445 0 0 $X=371850 $Y=184445
X928 1 MASCO__Y21 $T=371850 186445 0 0 $X=371850 $Y=186445
X929 1 MASCO__Y21 $T=371850 188445 0 0 $X=371850 $Y=188445
X930 1 MASCO__Y21 $T=379850 184445 0 0 $X=379850 $Y=184445
X931 1 MASCO__Y21 $T=379850 186445 0 0 $X=379850 $Y=186445
X932 1 MASCO__Y21 $T=379850 188445 0 0 $X=379850 $Y=188445
X933 1 MASCO__Y21 $T=387850 184445 0 0 $X=387850 $Y=184445
X934 1 MASCO__Y21 $T=387850 186445 0 0 $X=387850 $Y=186445
X935 1 MASCO__Y21 $T=387850 188445 0 0 $X=387850 $Y=188445
X936 1 MASCO__Y21 $T=395850 184445 0 0 $X=395850 $Y=184445
X937 1 MASCO__Y21 $T=395850 186445 0 0 $X=395850 $Y=186445
X938 1 MASCO__Y21 $T=395850 188445 0 0 $X=395850 $Y=188445
.ends MASCO__P5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: hvswitch5                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt hvswitch5 4 11 12 6 3 13 10 9 1
** N=13 EP=9 FDC=434
X0 1 2 3 4 MASCO__H1 $T=0 0 0 0 $X=251750 $Y=64655
X1 1 5 2 6 MASCO__H2 $T=0 0 0 0 $X=44775 $Y=96265
X2 1 7 8 6 2 MASCO__H3 $T=0 0 0 0 $X=84800 $Y=96265
X3 3 9 2 6 1 10 11 5 12 13
+ 7 4 MASCO__P4 $T=0 0 0 0 $X=-28920 $Y=-21375
X4 9 2 6 8 3 1 MASCO__P5 $T=0 0 0 0 $X=-28920 $Y=111955
.ends hvswitch5
