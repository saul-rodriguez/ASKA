* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : ref_bias                                     *
* Netlisted  : Mon Aug 26 08:30:34 2024                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(ne3) nem ndiff(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 1 MP(pe3) pem pdiff(D) p1trm(G) pdiff(S) nwtrm(B)
*.DEVTMPLT 2 NE3I_6() nemi_6 ndiff(D) p1trm(G) ndiff(S) pwitrm(B) dnwtrm(NW) bulk(SB)
*.DEVTMPLT 3 MOSVC3() mosvcm p1trm(G) nwtrm(NW) bulk(SB)
*.DEVTMPLT 4 D(p_dnw) p_dnw bulk(POS) nwtrm(NEG)
*.DEVTMPLT 5 D(p_ddnw) p_ddnw bulk(POS) dnwtrm(NEG)
*.DEVTMPLT 6 D(p_dipdnwmv) p_dipwmv pwitrm(POS) dnwtrm(NEG)
*.DEVTMPLT 7 D(p_dnw3) p_dnwm bulk(POS) nwtrm(NEG)
*.DEVTMPLT 8 R(rpp1k1_3) rpp1k1_s p1trm(POS) p1trm(NEG) bulk(SUB)
*.DEVTMPLT 9 C(cmm5t) cmim capm(POS) m4trm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_724653828770                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_724653828770 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_724653828770

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724653828771                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724653828771 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724653828771

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_724653828772                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_724653828772 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_724653828772

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724653828774                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724653828774 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724653828774

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724653828775                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724653828775 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724653828775

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724653828776                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724653828776 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724653828776

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724653828777                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724653828777 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724653828777

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724653828778                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724653828778 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724653828778

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724653828779                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724653828779 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724653828779

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246538287711                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246538287711 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246538287711

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246538287712                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246538287712 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246538287712

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246538287713                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246538287713 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246538287713

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246538287714                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246538287714 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246538287714

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246538287715                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246538287715 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246538287715

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246538287716                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246538287716 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246538287716

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246538287717                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246538287717 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246538287717

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246538287718                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246538287718 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246538287718

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246538287719                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246538287719 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246538287719

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246538287720                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246538287720 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246538287720

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246538287721                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246538287721 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246538287721

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_7246538287722                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_7246538287722 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_7246538287722

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246538287723                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246538287723 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246538287723

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246538287724                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246538287724 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246538287724

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246538287725                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246538287725 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246538287725

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246538287726                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246538287726 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246538287726

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246538287734                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246538287734 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246538287734

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246538287735                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246538287735 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7246538287735

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7246538287738                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7246538287738 1 2
** N=2 EP=2 FDC=0
.ends VIA1_C_CDNS_7246538287738

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724653828770                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724653828770 1 2 3 4 5
** N=5 EP=5 FDC=11
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=1
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=1
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=1
M4 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=6160 $Y=0 $dt=1
M5 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7700 $Y=0 $dt=1
M6 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=9240 $Y=0 $dt=1
M7 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10780 $Y=0 $dt=1
M8 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12320 $Y=0 $dt=1
M9 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=13860 $Y=0 $dt=1
D10 5 4 p_dnw3 AREA=2.15633e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=7
.ends pe3_CDNS_724653828770

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724653828771                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724653828771 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
.ends ne3_CDNS_724653828771

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724653828772                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724653828772 1 2 3 4 5
** N=5 EP=5 FDC=13
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=1
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=1
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=1
M4 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=6160 $Y=0 $dt=1
M5 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7700 $Y=0 $dt=1
M6 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=9240 $Y=0 $dt=1
M7 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10780 $Y=0 $dt=1
M8 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12320 $Y=0 $dt=1
M9 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=13860 $Y=0 $dt=1
M10 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=15400 $Y=0 $dt=1
M11 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=16940 $Y=0 $dt=1
D12 5 4 p_dnw3 AREA=2.52778e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=7
.ends pe3_CDNS_724653828772

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724653828773                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724653828773 1 2 3 4
** N=4 EP=4 FDC=3
M0 2 2 1 3 pe3 L=2e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 2 3 pe3 L=2e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=2540 $Y=0 $dt=1
D2 4 3 p_dnw3 AREA=9.11736e-11 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=7
.ends pe3_CDNS_724653828773

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_724653828774                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_724653828774 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.0005141 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=8
.ends rpp1k1_3_CDNS_724653828774

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724653828775                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724653828775 1 2 3 4
** N=4 EP=4 FDC=8
M0 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
M1 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=2540 $Y=0 $dt=0
M2 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=5080 $Y=0 $dt=0
M3 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7620 $Y=0 $dt=0
M4 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10160 $Y=0 $dt=0
M5 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12700 $Y=0 $dt=0
M6 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=15240 $Y=0 $dt=0
M7 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=17780 $Y=0 $dt=0
.ends ne3_CDNS_724653828775

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724653828779                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724653828779 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
M0 3 2 1 1 pe3 L=2e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_724653828779

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A1 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 2 3 6 pe3_CDNS_724653828779 $T=1510 1030 0 0 $X=0 $Y=0
X1 1 5 4 6 pe3_CDNS_724653828779 $T=4750 1030 0 0 $X=3240 $Y=0
.ends MASCO__A1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246538287710                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246538287710 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
M0 3 2 1 1 pe3 L=1e-05 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_7246538287710

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A2 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 4 2 6 pe3_CDNS_7246538287710 $T=1510 1030 0 0 $X=0 $Y=0
X1 1 5 3 6 pe3_CDNS_7246538287710 $T=12750 1030 0 0 $X=11240 $Y=0
.ends MASCO__A2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3i_6_CDNS_724653828778                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3i_6_CDNS_724653828778 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=1
X0 1 2 3 1 4 5 NE3I_6 w=1e-05 l=2e-06 as=4.8e-12 ad=4.8e-12 ps=2.096e-05 pd=2.096e-05 $X=0 $Y=0 $dt=2
.ends ne3i_6_CDNS_724653828778

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A3                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A3 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=2
X0 1 4 5 6 7 ne3i_6_CDNS_724653828778 $T=4060 14570 1 0 $X=0 $Y=0
X1 1 2 3 6 7 ne3i_6_CDNS_724653828778 $T=7460 14570 1 0 $X=3400 $Y=0
.ends MASCO__A3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A4                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A4 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=2
X0 1 4 5 6 7 ne3i_6_CDNS_724653828778 $T=4060 4450 0 0 $X=0 $Y=0
X1 1 2 3 6 7 ne3i_6_CDNS_724653828778 $T=7460 4450 0 0 $X=3400 $Y=0
.ends MASCO__A4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__B5                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__B5 1 2 3 4 5 6 7 8 9 10
+ 11
*.DEVICECLIMB
** N=11 EP=11 FDC=4
X0 1 10 6 5 3 2 11 MASCO__A3 $T=0 14680 0 0 $X=0 $Y=14680
X1 1 8 7 9 4 2 11 MASCO__A4 $T=0 0 0 0 $X=0 $Y=0
.ends MASCO__B5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A6                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A6 1 2 3 4 5 6 7 8
*.DEVICECLIMB
** N=8 EP=8 FDC=4
X0 1 2 3 5 4 8 MASCO__A1 $T=0 0 0 0 $X=0 $Y=0
X1 1 4 6 7 4 8 MASCO__A1 $T=6480 0 0 0 $X=6480 $Y=0
.ends MASCO__A6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ref_bias                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ref_bias 5 4 13 14 10 7 17
** N=18 EP=7 FDC=187
X0 1 VIA2_C_CDNS_724653828770 $T=13870 9200 0 0 $X=13160 $Y=8800
X1 1 VIA2_C_CDNS_724653828770 $T=13870 25290 0 0 $X=13160 $Y=24890
X2 2 VIA2_C_CDNS_724653828770 $T=64530 11760 0 0 $X=63820 $Y=11360
X3 2 VIA2_C_CDNS_724653828770 $T=64530 27850 0 0 $X=63820 $Y=27450
X4 3 VIA2_C_CDNS_724653828770 $T=66310 10480 0 0 $X=65600 $Y=10080
X5 3 VIA2_C_CDNS_724653828770 $T=66310 26570 0 0 $X=65600 $Y=26170
X6 4 VIA1_C_CDNS_724653828771 $T=17710 13040 0 0 $X=17570 $Y=12590
X7 4 VIA1_C_CDNS_724653828771 $T=17710 29130 0 0 $X=17570 $Y=28680
X8 4 VIA1_C_CDNS_724653828771 $T=20480 29130 0 0 $X=20340 $Y=28680
X9 4 VIA1_C_CDNS_724653828771 $T=20480 42300 0 0 $X=20340 $Y=41850
X10 4 VIA1_C_CDNS_724653828771 $T=23250 13040 0 0 $X=23110 $Y=12590
X11 4 VIA1_C_CDNS_724653828771 $T=23250 29130 0 0 $X=23110 $Y=28680
X12 4 VIA1_C_CDNS_724653828771 $T=23950 13040 0 0 $X=23810 $Y=12590
X13 4 VIA1_C_CDNS_724653828771 $T=23950 29130 0 0 $X=23810 $Y=28680
X14 1 VIA1_C_CDNS_724653828771 $T=26720 25290 0 0 $X=26580 $Y=24840
X15 3 VIA1_C_CDNS_724653828771 $T=29490 10480 0 0 $X=29350 $Y=10030
X16 1 VIA1_C_CDNS_724653828771 $T=29490 25290 0 0 $X=29350 $Y=24840
X17 4 VIA1_C_CDNS_724653828771 $T=30190 13040 0 0 $X=30050 $Y=12590
X18 4 VIA1_C_CDNS_724653828771 $T=30190 29130 0 0 $X=30050 $Y=28680
X19 1 VIA1_C_CDNS_724653828771 $T=32960 25290 0 0 $X=32820 $Y=24840
X20 1 VIA1_C_CDNS_724653828771 $T=35730 9200 0 0 $X=35590 $Y=8750
X21 3 VIA1_C_CDNS_724653828771 $T=35730 26570 0 0 $X=35590 $Y=26120
X22 4 VIA1_C_CDNS_724653828771 $T=36430 13040 0 0 $X=36290 $Y=12590
X23 4 VIA1_C_CDNS_724653828771 $T=36430 29130 0 0 $X=36290 $Y=28680
X24 1 VIA1_C_CDNS_724653828771 $T=39200 25290 0 0 $X=39060 $Y=24840
X25 2 VIA1_C_CDNS_724653828771 $T=41970 11760 0 0 $X=41830 $Y=11310
X26 1 VIA1_C_CDNS_724653828771 $T=41970 25290 0 0 $X=41830 $Y=24840
X27 4 VIA1_C_CDNS_724653828771 $T=42670 13040 0 0 $X=42530 $Y=12590
X28 4 VIA1_C_CDNS_724653828771 $T=42670 29130 0 0 $X=42530 $Y=28680
X29 1 VIA1_C_CDNS_724653828771 $T=45440 25290 0 0 $X=45300 $Y=24840
X30 1 VIA1_C_CDNS_724653828771 $T=48210 9200 0 0 $X=48070 $Y=8750
X31 3 VIA1_C_CDNS_724653828771 $T=48210 26570 0 0 $X=48070 $Y=26120
X32 4 VIA1_C_CDNS_724653828771 $T=48910 13040 0 0 $X=48770 $Y=12590
X33 4 VIA1_C_CDNS_724653828771 $T=48910 29130 0 0 $X=48770 $Y=28680
X34 1 VIA1_C_CDNS_724653828771 $T=51680 25290 0 0 $X=51540 $Y=24840
X35 4 VIA1_C_CDNS_724653828771 $T=51680 42300 0 0 $X=51540 $Y=41850
X36 3 VIA1_C_CDNS_724653828771 $T=54450 10480 0 0 $X=54310 $Y=10030
X37 4 VIA1_C_CDNS_724653828771 $T=54450 29130 0 0 $X=54310 $Y=28680
X38 4 VIA1_C_CDNS_724653828771 $T=55150 13040 0 0 $X=55010 $Y=12590
X39 4 VIA1_C_CDNS_724653828771 $T=55150 29130 0 0 $X=55010 $Y=28680
X40 4 VIA1_C_CDNS_724653828771 $T=57920 29130 0 0 $X=57780 $Y=28680
X41 4 VIA1_C_CDNS_724653828771 $T=57920 42300 0 0 $X=57780 $Y=41850
X42 4 VIA1_C_CDNS_724653828771 $T=60690 13040 0 0 $X=60550 $Y=12590
X43 4 VIA1_C_CDNS_724653828771 $T=60690 29130 0 0 $X=60550 $Y=28680
X44 4 VIA2_C_CDNS_724653828772 $T=15900 13040 0 0 $X=14930 $Y=12640
X45 4 VIA2_C_CDNS_724653828772 $T=15900 29130 0 0 $X=14930 $Y=28730
X46 4 VIA2_C_CDNS_724653828772 $T=15900 42300 0 0 $X=14930 $Y=41900
X47 4 VIA2_C_CDNS_724653828772 $T=62500 13040 0 0 $X=61530 $Y=12640
X48 4 VIA2_C_CDNS_724653828772 $T=62500 29130 0 0 $X=61530 $Y=28730
X49 4 VIA2_C_CDNS_724653828772 $T=62500 42300 0 0 $X=61530 $Y=41900
X50 1 VIA1_C_CDNS_724653828774 $T=26720 41270 0 0 $X=26580 $Y=41080
X51 1 VIA1_C_CDNS_724653828774 $T=32960 41270 0 0 $X=32820 $Y=41080
X52 1 VIA1_C_CDNS_724653828774 $T=39200 41270 0 0 $X=39060 $Y=41080
X53 1 VIA1_C_CDNS_724653828774 $T=45440 41270 0 0 $X=45300 $Y=41080
X54 1 VIA1_C_CDNS_724653828775 $T=17275 53125 0 0 $X=16875 $Y=52415
X55 5 VIA1_C_CDNS_724653828775 $T=19815 51345 0 0 $X=19415 $Y=50635
X56 1 VIA1_C_CDNS_724653828775 $T=22355 53125 0 0 $X=21955 $Y=52415
X57 5 VIA1_C_CDNS_724653828775 $T=24895 51345 0 0 $X=24495 $Y=50635
X58 1 VIA1_C_CDNS_724653828775 $T=27435 53125 0 0 $X=27035 $Y=52415
X59 5 VIA1_C_CDNS_724653828775 $T=29975 51345 0 0 $X=29575 $Y=50635
X60 1 VIA1_C_CDNS_724653828775 $T=32515 53125 0 0 $X=32115 $Y=52415
X61 5 VIA1_C_CDNS_724653828775 $T=35055 51345 0 0 $X=34655 $Y=50635
X62 1 VIA1_C_CDNS_724653828775 $T=37595 53125 0 0 $X=37195 $Y=52415
X63 3 VIA1_C_CDNS_724653828775 $T=42210 52905 0 0 $X=41810 $Y=52195
X64 6 VIA1_C_CDNS_724653828775 $T=44750 51125 0 0 $X=44350 $Y=50415
X65 3 VIA1_C_CDNS_724653828775 $T=47290 52905 0 0 $X=46890 $Y=52195
X66 6 VIA1_C_CDNS_724653828775 $T=49830 51125 0 0 $X=49430 $Y=50415
X67 3 VIA1_C_CDNS_724653828775 $T=52370 52905 0 0 $X=51970 $Y=52195
X68 6 VIA1_C_CDNS_724653828775 $T=54910 51125 0 0 $X=54510 $Y=50415
X69 3 VIA1_C_CDNS_724653828775 $T=57450 52905 0 0 $X=57050 $Y=52195
X70 6 VIA1_C_CDNS_724653828775 $T=59990 51125 0 0 $X=59590 $Y=50415
X71 3 VIA1_C_CDNS_724653828775 $T=62530 52905 0 0 $X=62130 $Y=52195
X72 7 VIA1_C_CDNS_724653828775 $T=137790 186425 0 0 $X=137390 $Y=185715
X73 8 VIA1_C_CDNS_724653828775 $T=140330 188205 0 0 $X=139930 $Y=187495
X74 7 VIA1_C_CDNS_724653828775 $T=142870 186425 0 0 $X=142470 $Y=185715
X75 8 VIA1_C_CDNS_724653828775 $T=147350 188205 0 0 $X=146950 $Y=187495
X76 2 VIA1_C_CDNS_724653828775 $T=149890 186425 0 0 $X=149490 $Y=185715
X77 8 VIA1_C_CDNS_724653828775 $T=152430 188205 0 0 $X=152030 $Y=187495
X78 9 VIA1_C_CDNS_724653828775 $T=162070 148400 0 0 $X=161670 $Y=147690
X79 10 VIA1_C_CDNS_724653828775 $T=163610 146620 0 0 $X=163210 $Y=145910
X80 9 VIA1_C_CDNS_724653828775 $T=165150 148400 0 0 $X=164750 $Y=147690
X81 7 VIA1_C_CDNS_724653828775 $T=165405 173875 0 0 $X=165005 $Y=173165
X82 7 VIA1_C_CDNS_724653828775 $T=165405 193895 0 0 $X=165005 $Y=193185
X83 7 VIA1_C_CDNS_724653828775 $T=166675 193895 0 0 $X=166275 $Y=193185
X84 7 VIA1_C_CDNS_724653828775 $T=166675 208575 0 0 $X=166275 $Y=207865
X85 10 VIA1_C_CDNS_724653828775 $T=166690 146620 0 0 $X=166290 $Y=145910
X86 7 VIA1_C_CDNS_724653828775 $T=167715 173875 0 0 $X=167315 $Y=173165
X87 7 VIA1_C_CDNS_724653828775 $T=167715 193895 0 0 $X=167315 $Y=193185
X88 9 VIA1_C_CDNS_724653828775 $T=168230 148400 0 0 $X=167830 $Y=147690
X89 7 VIA1_C_CDNS_724653828775 $T=168875 173875 0 0 $X=168475 $Y=173165
X90 7 VIA1_C_CDNS_724653828775 $T=168875 193895 0 0 $X=168475 $Y=193185
X91 10 VIA1_C_CDNS_724653828775 $T=169770 146620 0 0 $X=169370 $Y=145910
X92 11 VIA1_C_CDNS_724653828775 $T=170955 170315 0 0 $X=170555 $Y=169605
X93 12 VIA1_C_CDNS_724653828775 $T=170955 188555 0 0 $X=170555 $Y=187845
X94 9 VIA1_C_CDNS_724653828775 $T=171310 148400 0 0 $X=170910 $Y=147690
X95 7 VIA1_C_CDNS_724653828775 $T=172685 173875 0 0 $X=172285 $Y=173165
X96 7 VIA1_C_CDNS_724653828775 $T=172685 193895 0 0 $X=172285 $Y=193185
X97 10 VIA1_C_CDNS_724653828775 $T=172850 146620 0 0 $X=172450 $Y=145910
X98 12 VIA1_C_CDNS_724653828775 $T=174195 168535 0 0 $X=173795 $Y=167825
X99 9 VIA1_C_CDNS_724653828775 $T=174195 192115 0 0 $X=173795 $Y=191405
X100 9 VIA1_C_CDNS_724653828775 $T=174390 148400 0 0 $X=173990 $Y=147690
X101 7 VIA1_C_CDNS_724653828775 $T=175925 173875 0 0 $X=175525 $Y=173165
X102 7 VIA1_C_CDNS_724653828775 $T=175925 193895 0 0 $X=175525 $Y=193185
X103 10 VIA1_C_CDNS_724653828775 $T=175930 146620 0 0 $X=175530 $Y=145910
X104 9 VIA1_C_CDNS_724653828775 $T=177435 172095 0 0 $X=177035 $Y=171385
X105 11 VIA1_C_CDNS_724653828775 $T=177435 190335 0 0 $X=177035 $Y=189625
X106 9 VIA1_C_CDNS_724653828775 $T=177470 148400 0 0 $X=177070 $Y=147690
X107 10 VIA1_C_CDNS_724653828775 $T=179010 146620 0 0 $X=178610 $Y=145910
X108 7 VIA1_C_CDNS_724653828775 $T=179165 173875 0 0 $X=178765 $Y=173165
X109 7 VIA1_C_CDNS_724653828775 $T=179165 193895 0 0 $X=178765 $Y=193185
X110 9 VIA1_C_CDNS_724653828775 $T=180550 148400 0 0 $X=180150 $Y=147690
X111 11 VIA1_C_CDNS_724653828775 $T=180675 170315 0 0 $X=180275 $Y=169605
X112 12 VIA1_C_CDNS_724653828775 $T=180675 188555 0 0 $X=180275 $Y=187845
X113 7 VIA1_C_CDNS_724653828775 $T=182405 173875 0 0 $X=182005 $Y=173165
X114 7 VIA1_C_CDNS_724653828775 $T=182405 193895 0 0 $X=182005 $Y=193185
X115 9 VIA1_C_CDNS_724653828775 $T=183915 172095 0 0 $X=183515 $Y=171385
X116 12 VIA1_C_CDNS_724653828775 $T=183915 188555 0 0 $X=183515 $Y=187845
X117 7 VIA1_C_CDNS_724653828775 $T=185645 173875 0 0 $X=185245 $Y=173165
X118 7 VIA1_C_CDNS_724653828775 $T=185645 193895 0 0 $X=185245 $Y=193185
X119 12 VIA1_C_CDNS_724653828775 $T=187155 168535 0 0 $X=186755 $Y=167825
X120 9 VIA1_C_CDNS_724653828775 $T=187155 192115 0 0 $X=186755 $Y=191405
X121 7 VIA1_C_CDNS_724653828775 $T=188885 173875 0 0 $X=188485 $Y=173165
X122 7 VIA1_C_CDNS_724653828775 $T=188885 193895 0 0 $X=188485 $Y=193185
X123 11 VIA1_C_CDNS_724653828775 $T=189010 148400 0 0 $X=188610 $Y=147690
X124 9 VIA1_C_CDNS_724653828775 $T=190395 172095 0 0 $X=189995 $Y=171385
X125 11 VIA1_C_CDNS_724653828775 $T=190395 190335 0 0 $X=189995 $Y=189625
X126 13 VIA1_C_CDNS_724653828775 $T=190550 146620 0 0 $X=190150 $Y=145910
X127 11 VIA1_C_CDNS_724653828775 $T=192090 148400 0 0 $X=191690 $Y=147690
X128 7 VIA1_C_CDNS_724653828775 $T=192125 173875 0 0 $X=191725 $Y=173165
X129 7 VIA1_C_CDNS_724653828775 $T=192125 193895 0 0 $X=191725 $Y=193185
X130 13 VIA1_C_CDNS_724653828775 $T=193630 146620 0 0 $X=193230 $Y=145910
X131 11 VIA1_C_CDNS_724653828775 $T=193635 170315 0 0 $X=193235 $Y=169605
X132 9 VIA1_C_CDNS_724653828775 $T=193635 192115 0 0 $X=193235 $Y=191405
X133 11 VIA1_C_CDNS_724653828775 $T=195170 148400 0 0 $X=194770 $Y=147690
X134 7 VIA1_C_CDNS_724653828775 $T=195365 173875 0 0 $X=194965 $Y=173165
X135 7 VIA1_C_CDNS_724653828775 $T=195365 193895 0 0 $X=194965 $Y=193185
X136 13 VIA1_C_CDNS_724653828775 $T=196710 146620 0 0 $X=196310 $Y=145910
X137 9 VIA1_C_CDNS_724653828775 $T=196875 172095 0 0 $X=196475 $Y=171385
X138 12 VIA1_C_CDNS_724653828775 $T=196875 188555 0 0 $X=196475 $Y=187845
X139 11 VIA1_C_CDNS_724653828775 $T=198250 148400 0 0 $X=197850 $Y=147690
X140 7 VIA1_C_CDNS_724653828775 $T=198605 173875 0 0 $X=198205 $Y=173165
X141 7 VIA1_C_CDNS_724653828775 $T=198605 193895 0 0 $X=198205 $Y=193185
X142 13 VIA1_C_CDNS_724653828775 $T=199790 146620 0 0 $X=199390 $Y=145910
X143 12 VIA1_C_CDNS_724653828775 $T=200115 168535 0 0 $X=199715 $Y=167825
X144 9 VIA1_C_CDNS_724653828775 $T=200115 192115 0 0 $X=199715 $Y=191405
X145 11 VIA1_C_CDNS_724653828775 $T=201330 148400 0 0 $X=200930 $Y=147690
X146 7 VIA1_C_CDNS_724653828775 $T=201845 173875 0 0 $X=201445 $Y=173165
X147 7 VIA1_C_CDNS_724653828775 $T=201845 193895 0 0 $X=201445 $Y=193185
X148 13 VIA1_C_CDNS_724653828775 $T=202870 146620 0 0 $X=202470 $Y=145910
X149 9 VIA1_C_CDNS_724653828775 $T=203355 172095 0 0 $X=202955 $Y=171385
X150 11 VIA1_C_CDNS_724653828775 $T=203355 190335 0 0 $X=202955 $Y=189625
X151 11 VIA1_C_CDNS_724653828775 $T=204410 148400 0 0 $X=204010 $Y=147690
X152 7 VIA1_C_CDNS_724653828775 $T=205085 173875 0 0 $X=204685 $Y=173165
X153 7 VIA1_C_CDNS_724653828775 $T=205085 193895 0 0 $X=204685 $Y=193185
X154 11 VIA1_C_CDNS_724653828775 $T=206595 170315 0 0 $X=206195 $Y=169605
X155 9 VIA1_C_CDNS_724653828775 $T=206595 192115 0 0 $X=206195 $Y=191405
X156 7 VIA1_C_CDNS_724653828775 $T=208325 173875 0 0 $X=207925 $Y=173165
X157 7 VIA1_C_CDNS_724653828775 $T=208325 193895 0 0 $X=207925 $Y=193185
X158 11 VIA1_C_CDNS_724653828775 $T=209835 170315 0 0 $X=209435 $Y=169605
X159 12 VIA1_C_CDNS_724653828775 $T=209835 188555 0 0 $X=209435 $Y=187845
X160 7 VIA1_C_CDNS_724653828775 $T=211565 173875 0 0 $X=211165 $Y=173165
X161 7 VIA1_C_CDNS_724653828775 $T=211565 193895 0 0 $X=211165 $Y=193185
X162 12 VIA1_C_CDNS_724653828775 $T=212920 148400 0 0 $X=212520 $Y=147690
X163 12 VIA1_C_CDNS_724653828775 $T=213075 168535 0 0 $X=212675 $Y=167825
X164 9 VIA1_C_CDNS_724653828775 $T=213075 192115 0 0 $X=212675 $Y=191405
X165 14 VIA1_C_CDNS_724653828775 $T=214460 146620 0 0 $X=214060 $Y=145910
X166 7 VIA1_C_CDNS_724653828775 $T=214805 173875 0 0 $X=214405 $Y=173165
X167 7 VIA1_C_CDNS_724653828775 $T=214805 193895 0 0 $X=214405 $Y=193185
X168 12 VIA1_C_CDNS_724653828775 $T=216000 148400 0 0 $X=215600 $Y=147690
X169 9 VIA1_C_CDNS_724653828775 $T=216315 172095 0 0 $X=215915 $Y=171385
X170 11 VIA1_C_CDNS_724653828775 $T=216315 190335 0 0 $X=215915 $Y=189625
X171 14 VIA1_C_CDNS_724653828775 $T=217540 146620 0 0 $X=217140 $Y=145910
X172 7 VIA1_C_CDNS_724653828775 $T=218045 173875 0 0 $X=217645 $Y=173165
X173 7 VIA1_C_CDNS_724653828775 $T=218045 193895 0 0 $X=217645 $Y=193185
X174 12 VIA1_C_CDNS_724653828775 $T=219080 148400 0 0 $X=218680 $Y=147690
X175 11 VIA1_C_CDNS_724653828775 $T=219555 170315 0 0 $X=219155 $Y=169605
X176 12 VIA1_C_CDNS_724653828775 $T=219555 188555 0 0 $X=219155 $Y=187845
X177 14 VIA1_C_CDNS_724653828775 $T=220620 146620 0 0 $X=220220 $Y=145910
X178 7 VIA1_C_CDNS_724653828775 $T=221285 173875 0 0 $X=220885 $Y=173165
X179 7 VIA1_C_CDNS_724653828775 $T=221285 193895 0 0 $X=220885 $Y=193185
X180 7 VIA1_C_CDNS_724653828775 $T=221755 208575 0 0 $X=221355 $Y=207865
X181 12 VIA1_C_CDNS_724653828775 $T=222160 148400 0 0 $X=221760 $Y=147690
X182 7 VIA1_C_CDNS_724653828775 $T=223025 173875 0 0 $X=222625 $Y=173165
X183 7 VIA1_C_CDNS_724653828775 $T=223025 193895 0 0 $X=222625 $Y=193185
X184 14 VIA1_C_CDNS_724653828775 $T=223700 146620 0 0 $X=223300 $Y=145910
X185 12 VIA1_C_CDNS_724653828775 $T=225240 148400 0 0 $X=224840 $Y=147690
X186 14 VIA1_C_CDNS_724653828775 $T=226780 146620 0 0 $X=226380 $Y=145910
X187 12 VIA1_C_CDNS_724653828775 $T=228320 148400 0 0 $X=227920 $Y=147690
X188 2 VIA1_C_CDNS_724653828776 $T=162840 161880 0 0 $X=162440 $Y=161690
X189 2 VIA1_C_CDNS_724653828776 $T=164380 161880 0 0 $X=163980 $Y=161690
X190 2 VIA1_C_CDNS_724653828776 $T=165920 161880 0 0 $X=165520 $Y=161690
X191 2 VIA1_C_CDNS_724653828776 $T=167460 161880 0 0 $X=167060 $Y=161690
X192 2 VIA1_C_CDNS_724653828776 $T=169000 161880 0 0 $X=168600 $Y=161690
X193 2 VIA1_C_CDNS_724653828776 $T=170540 161880 0 0 $X=170140 $Y=161690
X194 2 VIA1_C_CDNS_724653828776 $T=172080 161880 0 0 $X=171680 $Y=161690
X195 2 VIA1_C_CDNS_724653828776 $T=173620 161880 0 0 $X=173220 $Y=161690
X196 2 VIA1_C_CDNS_724653828776 $T=175160 161880 0 0 $X=174760 $Y=161690
X197 2 VIA1_C_CDNS_724653828776 $T=176700 161880 0 0 $X=176300 $Y=161690
X198 2 VIA1_C_CDNS_724653828776 $T=178240 161880 0 0 $X=177840 $Y=161690
X199 2 VIA1_C_CDNS_724653828776 $T=179780 161880 0 0 $X=179380 $Y=161690
X200 2 VIA1_C_CDNS_724653828776 $T=189780 161880 0 0 $X=189380 $Y=161690
X201 2 VIA1_C_CDNS_724653828776 $T=191320 161880 0 0 $X=190920 $Y=161690
X202 2 VIA1_C_CDNS_724653828776 $T=192860 161880 0 0 $X=192460 $Y=161690
X203 2 VIA1_C_CDNS_724653828776 $T=194400 161880 0 0 $X=194000 $Y=161690
X204 2 VIA1_C_CDNS_724653828776 $T=195940 161880 0 0 $X=195540 $Y=161690
X205 2 VIA1_C_CDNS_724653828776 $T=197480 161880 0 0 $X=197080 $Y=161690
X206 2 VIA1_C_CDNS_724653828776 $T=199020 161880 0 0 $X=198620 $Y=161690
X207 2 VIA1_C_CDNS_724653828776 $T=200560 161880 0 0 $X=200160 $Y=161690
X208 2 VIA1_C_CDNS_724653828776 $T=202100 161880 0 0 $X=201700 $Y=161690
X209 2 VIA1_C_CDNS_724653828776 $T=203640 161880 0 0 $X=203240 $Y=161690
X210 2 VIA1_C_CDNS_724653828776 $T=213690 161880 0 0 $X=213290 $Y=161690
X211 2 VIA1_C_CDNS_724653828776 $T=215230 161880 0 0 $X=214830 $Y=161690
X212 2 VIA1_C_CDNS_724653828776 $T=216770 161880 0 0 $X=216370 $Y=161690
X213 2 VIA1_C_CDNS_724653828776 $T=218310 161880 0 0 $X=217910 $Y=161690
X214 2 VIA1_C_CDNS_724653828776 $T=219850 161880 0 0 $X=219450 $Y=161690
X215 2 VIA1_C_CDNS_724653828776 $T=221390 161880 0 0 $X=220990 $Y=161690
X216 2 VIA1_C_CDNS_724653828776 $T=222930 161880 0 0 $X=222530 $Y=161690
X217 2 VIA1_C_CDNS_724653828776 $T=224470 161880 0 0 $X=224070 $Y=161690
X218 2 VIA1_C_CDNS_724653828776 $T=226010 161880 0 0 $X=225610 $Y=161690
X219 2 VIA1_C_CDNS_724653828776 $T=227550 161880 0 0 $X=227150 $Y=161690
X220 5 VIA1_C_CDNS_724653828777 $T=18545 65405 0 0 $X=18355 $Y=65215
X221 5 VIA1_C_CDNS_724653828777 $T=21085 65405 0 0 $X=20895 $Y=65215
X222 5 VIA1_C_CDNS_724653828777 $T=23625 65405 0 0 $X=23435 $Y=65215
X223 5 VIA1_C_CDNS_724653828777 $T=26165 65405 0 0 $X=25975 $Y=65215
X224 5 VIA1_C_CDNS_724653828777 $T=28705 65405 0 0 $X=28515 $Y=65215
X225 5 VIA1_C_CDNS_724653828777 $T=31245 65405 0 0 $X=31055 $Y=65215
X226 5 VIA1_C_CDNS_724653828777 $T=33785 65405 0 0 $X=33595 $Y=65215
X227 5 VIA1_C_CDNS_724653828777 $T=36325 65405 0 0 $X=36135 $Y=65215
X228 5 VIA1_C_CDNS_724653828778 $T=43480 65295 0 0 $X=42560 $Y=65105
X229 5 VIA1_C_CDNS_724653828778 $T=46020 65295 0 0 $X=45100 $Y=65105
X230 5 VIA1_C_CDNS_724653828778 $T=48560 65295 0 0 $X=47640 $Y=65105
X231 5 VIA1_C_CDNS_724653828778 $T=51100 65295 0 0 $X=50180 $Y=65105
X232 5 VIA1_C_CDNS_724653828778 $T=53640 65295 0 0 $X=52720 $Y=65105
X233 5 VIA1_C_CDNS_724653828778 $T=56180 65295 0 0 $X=55260 $Y=65105
X234 5 VIA1_C_CDNS_724653828778 $T=58720 65295 0 0 $X=57800 $Y=65105
X235 5 VIA1_C_CDNS_724653828778 $T=61260 65295 0 0 $X=60340 $Y=65105
X236 8 VIA1_C_CDNS_724653828778 $T=139060 201685 0 0 $X=138140 $Y=201495
X237 8 VIA1_C_CDNS_724653828778 $T=141600 201685 0 0 $X=140680 $Y=201495
X238 2 VIA1_C_CDNS_724653828778 $T=148620 201685 0 0 $X=147700 $Y=201495
X239 2 VIA1_C_CDNS_724653828778 $T=151160 201685 0 0 $X=150240 $Y=201495
X240 7 VIA1_C_CDNS_724653828779 $T=22280 170260 0 0 $X=22140 $Y=169550
X241 7 VIA1_C_CDNS_724653828779 $T=22980 170260 0 0 $X=22840 $Y=169550
X242 7 VIA1_C_CDNS_724653828779 $T=22980 187940 0 0 $X=22840 $Y=187230
X243 15 VIA1_C_CDNS_724653828779 $T=33520 166700 0 0 $X=33380 $Y=165990
X244 16 VIA1_C_CDNS_724653828779 $T=33520 186160 0 0 $X=33380 $Y=185450
X245 7 VIA1_C_CDNS_724653828779 $T=34220 170260 0 0 $X=34080 $Y=169550
X246 7 VIA1_C_CDNS_724653828779 $T=34220 187940 0 0 $X=34080 $Y=187230
X247 16 VIA1_C_CDNS_724653828779 $T=44760 168480 0 0 $X=44620 $Y=167770
X248 15 VIA1_C_CDNS_724653828779 $T=44760 184380 0 0 $X=44620 $Y=183670
X249 7 VIA1_C_CDNS_724653828779 $T=45460 170260 0 0 $X=45320 $Y=169550
X250 7 VIA1_C_CDNS_724653828779 $T=45460 187940 0 0 $X=45320 $Y=187230
X251 15 VIA1_C_CDNS_724653828779 $T=56000 166700 0 0 $X=55860 $Y=165990
X252 16 VIA1_C_CDNS_724653828779 $T=56000 186160 0 0 $X=55860 $Y=185450
X253 7 VIA1_C_CDNS_724653828779 $T=56700 170260 0 0 $X=56560 $Y=169550
X254 7 VIA1_C_CDNS_724653828779 $T=56700 187940 0 0 $X=56560 $Y=187230
X255 16 VIA1_C_CDNS_724653828779 $T=67240 168480 0 0 $X=67100 $Y=167770
X256 15 VIA1_C_CDNS_724653828779 $T=67240 184380 0 0 $X=67100 $Y=183670
X257 7 VIA1_C_CDNS_724653828779 $T=67940 170260 0 0 $X=67800 $Y=169550
X258 7 VIA1_C_CDNS_724653828779 $T=67940 187940 0 0 $X=67800 $Y=187230
X259 15 VIA1_C_CDNS_724653828779 $T=78480 166700 0 0 $X=78340 $Y=165990
X260 16 VIA1_C_CDNS_724653828779 $T=78480 186160 0 0 $X=78340 $Y=185450
X261 7 VIA1_C_CDNS_724653828779 $T=79180 170260 0 0 $X=79040 $Y=169550
X262 7 VIA1_C_CDNS_724653828779 $T=79180 187940 0 0 $X=79040 $Y=187230
X263 16 VIA1_C_CDNS_724653828779 $T=89720 168480 0 0 $X=89580 $Y=167770
X264 15 VIA1_C_CDNS_724653828779 $T=89720 184380 0 0 $X=89580 $Y=183670
X265 7 VIA1_C_CDNS_724653828779 $T=90420 170260 0 0 $X=90280 $Y=169550
X266 7 VIA1_C_CDNS_724653828779 $T=90420 187940 0 0 $X=90280 $Y=187230
X267 15 VIA1_C_CDNS_724653828779 $T=100960 166700 0 0 $X=100820 $Y=165990
X268 16 VIA1_C_CDNS_724653828779 $T=100960 186160 0 0 $X=100820 $Y=185450
X269 7 VIA1_C_CDNS_724653828779 $T=101660 170260 0 0 $X=101520 $Y=169550
X270 7 VIA1_C_CDNS_724653828779 $T=101660 187940 0 0 $X=101520 $Y=187230
X271 16 VIA1_C_CDNS_724653828779 $T=112200 168480 0 0 $X=112060 $Y=167770
X272 15 VIA1_C_CDNS_724653828779 $T=112200 184380 0 0 $X=112060 $Y=183670
X273 7 VIA1_C_CDNS_724653828779 $T=112900 170260 0 0 $X=112760 $Y=169550
X274 7 VIA1_C_CDNS_724653828779 $T=112900 187940 0 0 $X=112760 $Y=187230
X275 15 VIA1_C_CDNS_7246538287711 $T=28250 201560 0 0 $X=27590 $Y=201370
X276 15 VIA1_C_CDNS_7246538287711 $T=39490 201560 0 0 $X=38830 $Y=201370
X277 15 VIA1_C_CDNS_7246538287711 $T=50730 201560 0 0 $X=50070 $Y=201370
X278 15 VIA1_C_CDNS_7246538287711 $T=61970 201560 0 0 $X=61310 $Y=201370
X279 15 VIA1_C_CDNS_7246538287711 $T=73210 201560 0 0 $X=72550 $Y=201370
X280 15 VIA1_C_CDNS_7246538287711 $T=84450 201560 0 0 $X=83790 $Y=201370
X281 15 VIA1_C_CDNS_7246538287711 $T=95690 201560 0 0 $X=95030 $Y=201370
X282 15 VIA1_C_CDNS_7246538287711 $T=106930 201560 0 0 $X=106270 $Y=201370
X283 16 VIA1_C_CDNS_7246538287712 $T=169915 187385 0 0 $X=168945 $Y=187195
X284 16 VIA1_C_CDNS_7246538287712 $T=169915 207405 0 0 $X=168945 $Y=207215
X285 16 VIA1_C_CDNS_7246538287712 $T=173155 187385 0 0 $X=172185 $Y=187195
X286 16 VIA1_C_CDNS_7246538287712 $T=173155 207405 0 0 $X=172185 $Y=207215
X287 16 VIA1_C_CDNS_7246538287712 $T=176395 187385 0 0 $X=175425 $Y=187195
X288 16 VIA1_C_CDNS_7246538287712 $T=176395 207405 0 0 $X=175425 $Y=207215
X289 16 VIA1_C_CDNS_7246538287712 $T=179635 187385 0 0 $X=178665 $Y=187195
X290 16 VIA1_C_CDNS_7246538287712 $T=179635 207405 0 0 $X=178665 $Y=207215
X291 16 VIA1_C_CDNS_7246538287712 $T=182875 187385 0 0 $X=181905 $Y=187195
X292 16 VIA1_C_CDNS_7246538287712 $T=182875 207405 0 0 $X=181905 $Y=207215
X293 16 VIA1_C_CDNS_7246538287712 $T=186115 187385 0 0 $X=185145 $Y=187195
X294 16 VIA1_C_CDNS_7246538287712 $T=186115 207405 0 0 $X=185145 $Y=207215
X295 16 VIA1_C_CDNS_7246538287712 $T=189355 187385 0 0 $X=188385 $Y=187195
X296 16 VIA1_C_CDNS_7246538287712 $T=189355 207405 0 0 $X=188385 $Y=207215
X297 16 VIA1_C_CDNS_7246538287712 $T=192595 187385 0 0 $X=191625 $Y=187195
X298 16 VIA1_C_CDNS_7246538287712 $T=192595 207405 0 0 $X=191625 $Y=207215
X299 16 VIA1_C_CDNS_7246538287712 $T=195835 187385 0 0 $X=194865 $Y=187195
X300 16 VIA1_C_CDNS_7246538287712 $T=195835 207405 0 0 $X=194865 $Y=207215
X301 16 VIA1_C_CDNS_7246538287712 $T=199075 187385 0 0 $X=198105 $Y=187195
X302 16 VIA1_C_CDNS_7246538287712 $T=199075 207405 0 0 $X=198105 $Y=207215
X303 16 VIA1_C_CDNS_7246538287712 $T=202315 187385 0 0 $X=201345 $Y=187195
X304 16 VIA1_C_CDNS_7246538287712 $T=202315 207405 0 0 $X=201345 $Y=207215
X305 16 VIA1_C_CDNS_7246538287712 $T=205555 187385 0 0 $X=204585 $Y=187195
X306 16 VIA1_C_CDNS_7246538287712 $T=205555 207405 0 0 $X=204585 $Y=207215
X307 16 VIA1_C_CDNS_7246538287712 $T=208795 187385 0 0 $X=207825 $Y=187195
X308 16 VIA1_C_CDNS_7246538287712 $T=208795 207405 0 0 $X=207825 $Y=207215
X309 16 VIA1_C_CDNS_7246538287712 $T=212035 187385 0 0 $X=211065 $Y=187195
X310 16 VIA1_C_CDNS_7246538287712 $T=212035 207405 0 0 $X=211065 $Y=207215
X311 16 VIA1_C_CDNS_7246538287712 $T=215275 187385 0 0 $X=214305 $Y=187195
X312 16 VIA1_C_CDNS_7246538287712 $T=215275 207405 0 0 $X=214305 $Y=207215
X313 16 VIA1_C_CDNS_7246538287712 $T=218515 187385 0 0 $X=217545 $Y=187195
X314 16 VIA1_C_CDNS_7246538287712 $T=218515 207405 0 0 $X=217545 $Y=207215
X315 7 VIA1_C_CDNS_7246538287713 $T=11740 170260 0 0 $X=11550 $Y=169600
X316 7 VIA1_C_CDNS_7246538287713 $T=11740 187940 0 0 $X=11550 $Y=187280
X317 7 VIA1_C_CDNS_7246538287713 $T=17010 187940 0 0 $X=16820 $Y=187280
X318 7 VIA1_C_CDNS_7246538287713 $T=22280 187940 0 0 $X=22090 $Y=187280
X319 15 VIA1_C_CDNS_7246538287713 $T=28250 184380 0 0 $X=28060 $Y=183720
X320 15 VIA1_C_CDNS_7246538287713 $T=39490 184380 0 0 $X=39300 $Y=183720
X321 15 VIA1_C_CDNS_7246538287713 $T=50730 184380 0 0 $X=50540 $Y=183720
X322 15 VIA1_C_CDNS_7246538287713 $T=61970 184380 0 0 $X=61780 $Y=183720
X323 15 VIA1_C_CDNS_7246538287713 $T=73210 184380 0 0 $X=73020 $Y=183720
X324 15 VIA1_C_CDNS_7246538287713 $T=84450 184380 0 0 $X=84260 $Y=183720
X325 15 VIA1_C_CDNS_7246538287713 $T=95690 184380 0 0 $X=95500 $Y=183720
X326 15 VIA1_C_CDNS_7246538287713 $T=106930 184380 0 0 $X=106740 $Y=183720
X327 7 VIA1_C_CDNS_7246538287713 $T=118170 187940 0 0 $X=117980 $Y=187280
X328 7 VIA1_C_CDNS_7246538287713 $T=123440 170260 0 0 $X=123250 $Y=169600
X329 7 VIA1_C_CDNS_7246538287713 $T=123440 187940 0 0 $X=123250 $Y=187280
X330 4 VIA2_C_CDNS_7246538287714 $T=15905 4500 0 0 $X=13335 $Y=3230
X331 4 VIA2_C_CDNS_7246538287714 $T=62500 4500 0 0 $X=59930 $Y=3230
X332 7 VIA2_C_CDNS_7246538287715 $T=9220 170260 0 0 $X=8250 $Y=169600
X333 7 VIA2_C_CDNS_7246538287715 $T=9220 187940 0 0 $X=8250 $Y=187280
X334 7 VIA2_C_CDNS_7246538287715 $T=125960 170260 0 0 $X=124990 $Y=169600
X335 7 VIA2_C_CDNS_7246538287715 $T=125960 187940 0 0 $X=124990 $Y=187280
X336 7 VIA2_C_CDNS_7246538287715 $T=162885 173875 0 0 $X=161915 $Y=173215
X337 7 VIA2_C_CDNS_7246538287715 $T=162885 193895 0 0 $X=161915 $Y=193235
X338 7 VIA2_C_CDNS_7246538287715 $T=162885 208575 0 0 $X=161915 $Y=207915
X339 7 VIA2_C_CDNS_7246538287715 $T=225545 173875 0 0 $X=224575 $Y=173215
X340 7 VIA2_C_CDNS_7246538287715 $T=225545 193895 0 0 $X=224575 $Y=193235
X341 7 VIA2_C_CDNS_7246538287715 $T=225545 208575 0 0 $X=224575 $Y=207915
X342 15 VIA2_C_CDNS_7246538287716 $T=7190 166700 0 0 $X=6480 $Y=166040
X343 15 VIA2_C_CDNS_7246538287716 $T=7190 184380 0 0 $X=6480 $Y=183720
X344 16 VIA2_C_CDNS_7246538287716 $T=127990 168480 0 0 $X=127280 $Y=167820
X345 16 VIA2_C_CDNS_7246538287716 $T=127990 186160 0 0 $X=127280 $Y=185500
X346 9 VIA2_C_CDNS_7246538287716 $T=160855 172095 0 0 $X=160145 $Y=171435
X347 9 VIA2_C_CDNS_7246538287716 $T=160855 192115 0 0 $X=160145 $Y=191455
X348 11 VIA2_C_CDNS_7246538287716 $T=227575 170315 0 0 $X=226865 $Y=169655
X349 11 VIA2_C_CDNS_7246538287716 $T=227575 190335 0 0 $X=226865 $Y=189675
X350 12 VIA2_C_CDNS_7246538287716 $T=229355 168535 0 0 $X=228645 $Y=167875
X351 12 VIA2_C_CDNS_7246538287716 $T=229355 188555 0 0 $X=228645 $Y=187895
X352 4 VIA1_C_CDNS_7246538287717 $T=117240 7840 0 90 $X=116270 $Y=7440
X353 4 VIA1_C_CDNS_7246538287717 $T=117240 38150 0 90 $X=116270 $Y=37750
X354 4 VIA1_C_CDNS_7246538287717 $T=117240 39310 0 90 $X=116270 $Y=38910
X355 4 VIA1_C_CDNS_7246538287717 $T=117240 69390 0 90 $X=116270 $Y=68990
X356 4 VIA1_C_CDNS_7246538287717 $T=117240 70550 0 90 $X=116270 $Y=70150
X357 4 VIA1_C_CDNS_7246538287717 $T=117240 100860 0 90 $X=116270 $Y=100460
X358 4 VIA1_C_CDNS_7246538287717 $T=154205 7780 0 90 $X=153235 $Y=7380
X359 4 VIA1_C_CDNS_7246538287717 $T=154205 38090 0 90 $X=153235 $Y=37690
X360 4 VIA1_C_CDNS_7246538287717 $T=154205 39250 0 90 $X=153235 $Y=38850
X361 4 VIA1_C_CDNS_7246538287717 $T=154205 69330 0 90 $X=153235 $Y=68930
X362 4 VIA1_C_CDNS_7246538287717 $T=154205 70490 0 90 $X=153235 $Y=70090
X363 4 VIA1_C_CDNS_7246538287717 $T=154205 100800 0 90 $X=153235 $Y=100400
X364 14 VIA1_C_CDNS_7246538287718 $T=83930 23110 0 90 $X=83220 $Y=22450
X365 14 VIA1_C_CDNS_7246538287718 $T=83930 54350 0 90 $X=83220 $Y=53690
X366 14 VIA1_C_CDNS_7246538287718 $T=83930 85590 0 90 $X=83220 $Y=84930
X367 13 VIA1_C_CDNS_7246538287718 $T=120895 23050 0 90 $X=120185 $Y=22390
X368 13 VIA1_C_CDNS_7246538287718 $T=120895 54290 0 90 $X=120185 $Y=53630
X369 13 VIA1_C_CDNS_7246538287718 $T=120895 85530 0 90 $X=120185 $Y=84870
X370 10 VIA2_C_CDNS_7246538287719 $T=17790 130490 0 0 $X=17650 $Y=130300
X371 17 VIA2_C_CDNS_7246538287719 $T=17790 131270 0 0 $X=17650 $Y=131080
X372 10 VIA2_C_CDNS_7246538287719 $T=20880 130490 0 0 $X=20740 $Y=130300
X373 17 VIA2_C_CDNS_7246538287719 $T=21500 131270 0 0 $X=21360 $Y=131080
X374 10 VIA2_C_CDNS_7246538287719 $T=24590 130490 0 0 $X=24450 $Y=130300
X375 17 VIA2_C_CDNS_7246538287719 $T=24590 131270 0 0 $X=24450 $Y=131080
X376 10 VIA2_C_CDNS_7246538287719 $T=27680 130490 0 0 $X=27540 $Y=130300
X377 17 VIA2_C_CDNS_7246538287719 $T=28300 131270 0 0 $X=28160 $Y=131080
X378 10 VIA2_C_CDNS_7246538287719 $T=31390 130490 0 0 $X=31250 $Y=130300
X379 17 VIA2_C_CDNS_7246538287719 $T=31390 131270 0 0 $X=31250 $Y=131080
X380 10 VIA2_C_CDNS_7246538287719 $T=34480 130490 0 0 $X=34340 $Y=130300
X381 17 VIA2_C_CDNS_7246538287719 $T=35100 131270 0 0 $X=34960 $Y=131080
X382 10 VIA2_C_CDNS_7246538287719 $T=38190 130490 0 0 $X=38050 $Y=130300
X383 17 VIA2_C_CDNS_7246538287719 $T=38190 131270 0 0 $X=38050 $Y=131080
X384 10 VIA2_C_CDNS_7246538287719 $T=41280 130490 0 0 $X=41140 $Y=130300
X385 17 VIA2_C_CDNS_7246538287719 $T=41900 131270 0 0 $X=41760 $Y=131080
X386 10 VIA2_C_CDNS_7246538287719 $T=44990 130490 0 0 $X=44850 $Y=130300
X387 17 VIA2_C_CDNS_7246538287719 $T=44990 131270 0 0 $X=44850 $Y=131080
X388 10 VIA2_C_CDNS_7246538287719 $T=48080 130490 0 0 $X=47940 $Y=130300
X389 17 VIA2_C_CDNS_7246538287719 $T=48700 131270 0 0 $X=48560 $Y=131080
X390 10 VIA2_C_CDNS_7246538287719 $T=51790 130490 0 0 $X=51650 $Y=130300
X391 17 VIA2_C_CDNS_7246538287719 $T=51790 131270 0 0 $X=51650 $Y=131080
X392 10 VIA2_C_CDNS_7246538287719 $T=54880 130490 0 0 $X=54740 $Y=130300
X393 17 VIA2_C_CDNS_7246538287719 $T=55500 131270 0 0 $X=55360 $Y=131080
X394 10 VIA2_C_CDNS_7246538287719 $T=58590 130490 0 0 $X=58450 $Y=130300
X395 17 VIA2_C_CDNS_7246538287719 $T=58590 131270 0 0 $X=58450 $Y=131080
X396 10 VIA2_C_CDNS_7246538287719 $T=61680 130490 0 0 $X=61540 $Y=130300
X397 17 VIA2_C_CDNS_7246538287719 $T=62300 131270 0 0 $X=62160 $Y=131080
X398 6 VIA1_C_CDNS_7246538287720 $T=14390 117740 0 0 $X=13680 $Y=117600
X399 6 VIA1_C_CDNS_7246538287720 $T=14390 144020 0 0 $X=13680 $Y=143880
X400 6 VIA1_C_CDNS_7246538287720 $T=17790 117740 0 0 $X=17080 $Y=117600
X401 6 VIA1_C_CDNS_7246538287720 $T=17790 144020 0 0 $X=17080 $Y=143880
X402 6 VIA1_C_CDNS_7246538287720 $T=21190 117740 0 0 $X=20480 $Y=117600
X403 6 VIA1_C_CDNS_7246538287720 $T=21190 144020 0 0 $X=20480 $Y=143880
X404 6 VIA1_C_CDNS_7246538287720 $T=24590 117740 0 0 $X=23880 $Y=117600
X405 6 VIA1_C_CDNS_7246538287720 $T=24590 144020 0 0 $X=23880 $Y=143880
X406 6 VIA1_C_CDNS_7246538287720 $T=27990 117740 0 0 $X=27280 $Y=117600
X407 6 VIA1_C_CDNS_7246538287720 $T=27990 144020 0 0 $X=27280 $Y=143880
X408 6 VIA1_C_CDNS_7246538287720 $T=31390 117740 0 0 $X=30680 $Y=117600
X409 6 VIA1_C_CDNS_7246538287720 $T=31390 144020 0 0 $X=30680 $Y=143880
X410 6 VIA1_C_CDNS_7246538287720 $T=34790 117740 0 0 $X=34080 $Y=117600
X411 6 VIA1_C_CDNS_7246538287720 $T=34790 144020 0 0 $X=34080 $Y=143880
X412 6 VIA1_C_CDNS_7246538287720 $T=38190 117740 0 0 $X=37480 $Y=117600
X413 6 VIA1_C_CDNS_7246538287720 $T=38190 144020 0 0 $X=37480 $Y=143880
X414 6 VIA1_C_CDNS_7246538287720 $T=41590 117740 0 0 $X=40880 $Y=117600
X415 6 VIA1_C_CDNS_7246538287720 $T=41590 144020 0 0 $X=40880 $Y=143880
X416 6 VIA1_C_CDNS_7246538287720 $T=44990 117740 0 0 $X=44280 $Y=117600
X417 6 VIA1_C_CDNS_7246538287720 $T=44990 144020 0 0 $X=44280 $Y=143880
X418 6 VIA1_C_CDNS_7246538287720 $T=48390 117740 0 0 $X=47680 $Y=117600
X419 6 VIA1_C_CDNS_7246538287720 $T=48390 144020 0 0 $X=47680 $Y=143880
X420 6 VIA1_C_CDNS_7246538287720 $T=51790 117740 0 0 $X=51080 $Y=117600
X421 6 VIA1_C_CDNS_7246538287720 $T=51790 144020 0 0 $X=51080 $Y=143880
X422 6 VIA1_C_CDNS_7246538287720 $T=55190 117740 0 0 $X=54480 $Y=117600
X423 6 VIA1_C_CDNS_7246538287720 $T=55190 144020 0 0 $X=54480 $Y=143880
X424 6 VIA1_C_CDNS_7246538287720 $T=58590 117740 0 0 $X=57880 $Y=117600
X425 6 VIA1_C_CDNS_7246538287720 $T=58590 144020 0 0 $X=57880 $Y=143880
X426 6 VIA1_C_CDNS_7246538287720 $T=61990 117740 0 0 $X=61280 $Y=117600
X427 6 VIA1_C_CDNS_7246538287720 $T=61990 144020 0 0 $X=61280 $Y=143880
X428 6 VIA1_C_CDNS_7246538287720 $T=65390 117740 0 0 $X=64680 $Y=117600
X429 6 VIA1_C_CDNS_7246538287720 $T=65390 144020 0 0 $X=64680 $Y=143880
X430 6 VIA2_C_CDNS_7246538287721 $T=13120 115960 0 0 $X=12980 $Y=115250
X431 6 VIA2_C_CDNS_7246538287721 $T=13120 145800 0 0 $X=12980 $Y=145090
X432 6 VIA2_C_CDNS_7246538287721 $T=14390 115960 0 0 $X=14250 $Y=115250
X433 6 VIA2_C_CDNS_7246538287721 $T=14390 145800 0 0 $X=14250 $Y=145090
X434 6 VIA2_C_CDNS_7246538287721 $T=15660 115960 0 0 $X=15520 $Y=115250
X435 6 VIA2_C_CDNS_7246538287721 $T=15660 145800 0 0 $X=15520 $Y=145090
X436 6 VIA2_C_CDNS_7246538287721 $T=16520 115960 0 0 $X=16380 $Y=115250
X437 6 VIA2_C_CDNS_7246538287721 $T=16520 145800 0 0 $X=16380 $Y=145090
X438 6 VIA2_C_CDNS_7246538287721 $T=17790 115960 0 0 $X=17650 $Y=115250
X439 6 VIA2_C_CDNS_7246538287721 $T=17790 145800 0 0 $X=17650 $Y=145090
X440 15 VIA2_C_CDNS_7246538287721 $T=19060 112400 0 0 $X=18920 $Y=111690
X441 16 VIA2_C_CDNS_7246538287721 $T=19060 149360 0 0 $X=18920 $Y=148650
X442 6 VIA2_C_CDNS_7246538287721 $T=19920 115960 0 0 $X=19780 $Y=115250
X443 6 VIA2_C_CDNS_7246538287721 $T=19920 145800 0 0 $X=19780 $Y=145090
X444 6 VIA2_C_CDNS_7246538287721 $T=21190 115960 0 0 $X=21050 $Y=115250
X445 6 VIA2_C_CDNS_7246538287721 $T=21190 145800 0 0 $X=21050 $Y=145090
X446 16 VIA2_C_CDNS_7246538287721 $T=22460 114180 0 0 $X=22320 $Y=113470
X447 15 VIA2_C_CDNS_7246538287721 $T=22460 147580 0 0 $X=22320 $Y=146870
X448 6 VIA2_C_CDNS_7246538287721 $T=23320 115960 0 0 $X=23180 $Y=115250
X449 6 VIA2_C_CDNS_7246538287721 $T=23320 145800 0 0 $X=23180 $Y=145090
X450 6 VIA2_C_CDNS_7246538287721 $T=24590 115960 0 0 $X=24450 $Y=115250
X451 6 VIA2_C_CDNS_7246538287721 $T=24590 145800 0 0 $X=24450 $Y=145090
X452 15 VIA2_C_CDNS_7246538287721 $T=25860 112400 0 0 $X=25720 $Y=111690
X453 16 VIA2_C_CDNS_7246538287721 $T=25860 149360 0 0 $X=25720 $Y=148650
X454 6 VIA2_C_CDNS_7246538287721 $T=26720 115960 0 0 $X=26580 $Y=115250
X455 6 VIA2_C_CDNS_7246538287721 $T=26720 145800 0 0 $X=26580 $Y=145090
X456 6 VIA2_C_CDNS_7246538287721 $T=27990 115960 0 0 $X=27850 $Y=115250
X457 6 VIA2_C_CDNS_7246538287721 $T=27990 145800 0 0 $X=27850 $Y=145090
X458 16 VIA2_C_CDNS_7246538287721 $T=29260 114180 0 0 $X=29120 $Y=113470
X459 15 VIA2_C_CDNS_7246538287721 $T=29260 147580 0 0 $X=29120 $Y=146870
X460 6 VIA2_C_CDNS_7246538287721 $T=30120 115960 0 0 $X=29980 $Y=115250
X461 6 VIA2_C_CDNS_7246538287721 $T=30120 145800 0 0 $X=29980 $Y=145090
X462 6 VIA2_C_CDNS_7246538287721 $T=31390 115960 0 0 $X=31250 $Y=115250
X463 6 VIA2_C_CDNS_7246538287721 $T=31390 145800 0 0 $X=31250 $Y=145090
X464 15 VIA2_C_CDNS_7246538287721 $T=32660 112400 0 0 $X=32520 $Y=111690
X465 16 VIA2_C_CDNS_7246538287721 $T=32660 149360 0 0 $X=32520 $Y=148650
X466 6 VIA2_C_CDNS_7246538287721 $T=33520 115960 0 0 $X=33380 $Y=115250
X467 6 VIA2_C_CDNS_7246538287721 $T=33520 145800 0 0 $X=33380 $Y=145090
X468 6 VIA2_C_CDNS_7246538287721 $T=34790 115960 0 0 $X=34650 $Y=115250
X469 6 VIA2_C_CDNS_7246538287721 $T=34790 145800 0 0 $X=34650 $Y=145090
X470 16 VIA2_C_CDNS_7246538287721 $T=36060 114180 0 0 $X=35920 $Y=113470
X471 15 VIA2_C_CDNS_7246538287721 $T=36060 147580 0 0 $X=35920 $Y=146870
X472 6 VIA2_C_CDNS_7246538287721 $T=36920 115960 0 0 $X=36780 $Y=115250
X473 6 VIA2_C_CDNS_7246538287721 $T=36920 145800 0 0 $X=36780 $Y=145090
X474 6 VIA2_C_CDNS_7246538287721 $T=38190 115960 0 0 $X=38050 $Y=115250
X475 6 VIA2_C_CDNS_7246538287721 $T=38190 145800 0 0 $X=38050 $Y=145090
X476 15 VIA2_C_CDNS_7246538287721 $T=39460 112400 0 0 $X=39320 $Y=111690
X477 16 VIA2_C_CDNS_7246538287721 $T=39460 149360 0 0 $X=39320 $Y=148650
X478 6 VIA2_C_CDNS_7246538287721 $T=40320 115960 0 0 $X=40180 $Y=115250
X479 6 VIA2_C_CDNS_7246538287721 $T=40320 145800 0 0 $X=40180 $Y=145090
X480 6 VIA2_C_CDNS_7246538287721 $T=41590 115960 0 0 $X=41450 $Y=115250
X481 6 VIA2_C_CDNS_7246538287721 $T=41590 145800 0 0 $X=41450 $Y=145090
X482 16 VIA2_C_CDNS_7246538287721 $T=42860 114180 0 0 $X=42720 $Y=113470
X483 15 VIA2_C_CDNS_7246538287721 $T=42860 147580 0 0 $X=42720 $Y=146870
X484 6 VIA2_C_CDNS_7246538287721 $T=43720 115960 0 0 $X=43580 $Y=115250
X485 6 VIA2_C_CDNS_7246538287721 $T=43720 145800 0 0 $X=43580 $Y=145090
X486 6 VIA2_C_CDNS_7246538287721 $T=44990 115960 0 0 $X=44850 $Y=115250
X487 6 VIA2_C_CDNS_7246538287721 $T=44990 145800 0 0 $X=44850 $Y=145090
X488 15 VIA2_C_CDNS_7246538287721 $T=46260 112400 0 0 $X=46120 $Y=111690
X489 16 VIA2_C_CDNS_7246538287721 $T=46260 149360 0 0 $X=46120 $Y=148650
X490 6 VIA2_C_CDNS_7246538287721 $T=47120 115960 0 0 $X=46980 $Y=115250
X491 6 VIA2_C_CDNS_7246538287721 $T=47120 145800 0 0 $X=46980 $Y=145090
X492 6 VIA2_C_CDNS_7246538287721 $T=48390 115960 0 0 $X=48250 $Y=115250
X493 6 VIA2_C_CDNS_7246538287721 $T=48390 145800 0 0 $X=48250 $Y=145090
X494 16 VIA2_C_CDNS_7246538287721 $T=49660 114180 0 0 $X=49520 $Y=113470
X495 15 VIA2_C_CDNS_7246538287721 $T=49660 147580 0 0 $X=49520 $Y=146870
X496 6 VIA2_C_CDNS_7246538287721 $T=50520 115960 0 0 $X=50380 $Y=115250
X497 6 VIA2_C_CDNS_7246538287721 $T=50520 145800 0 0 $X=50380 $Y=145090
X498 6 VIA2_C_CDNS_7246538287721 $T=51790 115960 0 0 $X=51650 $Y=115250
X499 6 VIA2_C_CDNS_7246538287721 $T=51790 145800 0 0 $X=51650 $Y=145090
X500 15 VIA2_C_CDNS_7246538287721 $T=53060 112400 0 0 $X=52920 $Y=111690
X501 16 VIA2_C_CDNS_7246538287721 $T=53060 149360 0 0 $X=52920 $Y=148650
X502 6 VIA2_C_CDNS_7246538287721 $T=53920 115960 0 0 $X=53780 $Y=115250
X503 6 VIA2_C_CDNS_7246538287721 $T=53920 145800 0 0 $X=53780 $Y=145090
X504 6 VIA2_C_CDNS_7246538287721 $T=55190 115960 0 0 $X=55050 $Y=115250
X505 6 VIA2_C_CDNS_7246538287721 $T=55190 145800 0 0 $X=55050 $Y=145090
X506 16 VIA2_C_CDNS_7246538287721 $T=56460 114180 0 0 $X=56320 $Y=113470
X507 15 VIA2_C_CDNS_7246538287721 $T=56460 147580 0 0 $X=56320 $Y=146870
X508 6 VIA2_C_CDNS_7246538287721 $T=57320 115960 0 0 $X=57180 $Y=115250
X509 6 VIA2_C_CDNS_7246538287721 $T=57320 145800 0 0 $X=57180 $Y=145090
X510 6 VIA2_C_CDNS_7246538287721 $T=58590 115960 0 0 $X=58450 $Y=115250
X511 6 VIA2_C_CDNS_7246538287721 $T=58590 145800 0 0 $X=58450 $Y=145090
X512 15 VIA2_C_CDNS_7246538287721 $T=59860 112400 0 0 $X=59720 $Y=111690
X513 16 VIA2_C_CDNS_7246538287721 $T=59860 149360 0 0 $X=59720 $Y=148650
X514 6 VIA2_C_CDNS_7246538287721 $T=60720 115960 0 0 $X=60580 $Y=115250
X515 6 VIA2_C_CDNS_7246538287721 $T=60720 145800 0 0 $X=60580 $Y=145090
X516 6 VIA2_C_CDNS_7246538287721 $T=61990 115960 0 0 $X=61850 $Y=115250
X517 6 VIA2_C_CDNS_7246538287721 $T=61990 145800 0 0 $X=61850 $Y=145090
X518 16 VIA2_C_CDNS_7246538287721 $T=63260 114180 0 0 $X=63120 $Y=113470
X519 15 VIA2_C_CDNS_7246538287721 $T=63260 147580 0 0 $X=63120 $Y=146870
X520 6 VIA2_C_CDNS_7246538287721 $T=64120 115960 0 0 $X=63980 $Y=115250
X521 6 VIA2_C_CDNS_7246538287721 $T=64120 145800 0 0 $X=63980 $Y=145090
X522 6 VIA2_C_CDNS_7246538287721 $T=65390 115960 0 0 $X=65250 $Y=115250
X523 6 VIA2_C_CDNS_7246538287721 $T=65390 145800 0 0 $X=65250 $Y=145090
X524 6 VIA2_C_CDNS_7246538287721 $T=66660 115960 0 0 $X=66520 $Y=115250
X525 6 VIA2_C_CDNS_7246538287721 $T=66660 145800 0 0 $X=66520 $Y=145090
X526 15 VIA3_C_CDNS_7246538287722 $T=7620 112400 0 0 $X=6910 $Y=111740
X527 15 VIA3_C_CDNS_7246538287722 $T=7620 147580 0 0 $X=6910 $Y=146920
X528 16 VIA3_C_CDNS_7246538287722 $T=9500 114180 0 0 $X=8790 $Y=113520
X529 16 VIA3_C_CDNS_7246538287722 $T=9500 149360 0 0 $X=8790 $Y=148700
X530 6 VIA3_C_CDNS_7246538287722 $T=11380 115960 0 0 $X=10670 $Y=115300
X531 6 VIA3_C_CDNS_7246538287722 $T=11380 145800 0 0 $X=10670 $Y=145140
X532 6 VIA3_C_CDNS_7246538287722 $T=68400 115960 0 0 $X=67690 $Y=115300
X533 6 VIA3_C_CDNS_7246538287722 $T=68400 145800 0 0 $X=67690 $Y=145140
X534 15 VIA3_C_CDNS_7246538287722 $T=70280 112400 0 0 $X=69570 $Y=111740
X535 15 VIA3_C_CDNS_7246538287722 $T=70280 147580 0 0 $X=69570 $Y=146920
X536 16 VIA3_C_CDNS_7246538287722 $T=72160 114180 0 0 $X=71450 $Y=113520
X537 16 VIA3_C_CDNS_7246538287722 $T=72160 149360 0 0 $X=71450 $Y=148700
X538 4 VIA1_C_CDNS_7246538287723 $T=15905 4500 0 0 $X=13335 $Y=3230
X539 4 VIA1_C_CDNS_7246538287723 $T=62500 4500 0 0 $X=59930 $Y=3230
X540 1 VIA2_C_CDNS_7246538287724 $T=17575 53125 0 0 $X=16825 $Y=52375
X541 9 VIA2_C_CDNS_7246538287724 $T=163125 148400 0 0 $X=162375 $Y=147650
X542 11 VIA2_C_CDNS_7246538287724 $T=204535 148400 0 0 $X=203785 $Y=147650
X543 12 VIA2_C_CDNS_7246538287724 $T=226740 148400 0 0 $X=225990 $Y=147650
X544 2 VIA2_C_CDNS_7246538287725 $T=152805 186425 0 0 $X=152055 $Y=185675
X545 14 VIA2_C_CDNS_7246538287725 $T=187300 141530 0 0 $X=186550 $Y=140780
X546 10 VIA2_C_CDNS_7246538287726 $T=170630 146620 0 0 $X=168580 $Y=145870
X547 13 VIA2_C_CDNS_7246538287726 $T=196715 146620 0 0 $X=194665 $Y=145870
X548 14 VIA2_C_CDNS_7246538287726 $T=220620 146620 0 0 $X=218570 $Y=145870
X549 18 VIA2_C_CDNS_7246538287734 $T=82800 119325 0 0 $X=82310 $Y=117275
X550 10 VIA2_C_CDNS_7246538287734 $T=82850 149150 0 0 $X=82360 $Y=147100
X551 18 VIA1_C_CDNS_7246538287735 $T=82800 119325 0 0 $X=82310 $Y=117275
X552 10 VIA1_C_CDNS_7246538287735 $T=82850 149150 0 0 $X=82360 $Y=147100
X553 7 4 VIA1_C_CDNS_7246538287738 $T=70935 208110 0 0 $X=65765 $Y=205540
X554 7 4 VIA1_C_CDNS_7246538287738 $T=150700 208200 0 0 $X=145530 $Y=205630
X555 11 2 13 7 4 pe3_CDNS_724653828770 $T=189280 150320 0 0 $X=187770 $Y=149290
X556 12 2 14 7 4 pe3_CDNS_724653828770 $T=213190 150320 0 0 $X=211680 $Y=149290
X557 4 4 4 ne3_CDNS_724653828771 $T=17980 14080 0 0 $X=17180 $Y=13680
X558 4 4 4 ne3_CDNS_724653828771 $T=17980 30170 0 0 $X=17180 $Y=29770
X559 4 1 3 ne3_CDNS_724653828771 $T=24220 14080 0 0 $X=23420 $Y=13680
X560 4 1 1 ne3_CDNS_724653828771 $T=24220 30170 0 0 $X=23420 $Y=29770
X561 4 1 1 ne3_CDNS_724653828771 $T=30460 14080 0 0 $X=29660 $Y=13680
X562 4 1 3 ne3_CDNS_724653828771 $T=30460 30170 0 0 $X=29660 $Y=29770
X563 4 1 2 ne3_CDNS_724653828771 $T=36700 14080 0 0 $X=35900 $Y=13680
X564 4 1 1 ne3_CDNS_724653828771 $T=36700 30170 0 0 $X=35900 $Y=29770
X565 4 1 1 ne3_CDNS_724653828771 $T=42940 14080 0 0 $X=42140 $Y=13680
X566 4 1 3 ne3_CDNS_724653828771 $T=42940 30170 0 0 $X=42140 $Y=29770
X567 4 1 3 ne3_CDNS_724653828771 $T=49180 14080 0 0 $X=48380 $Y=13680
X568 4 4 4 ne3_CDNS_724653828771 $T=49180 30170 0 0 $X=48380 $Y=29770
X569 4 4 4 ne3_CDNS_724653828771 $T=55420 14080 0 0 $X=54620 $Y=13680
X570 4 4 4 ne3_CDNS_724653828771 $T=55420 30170 0 0 $X=54620 $Y=29770
X571 9 2 10 7 4 pe3_CDNS_724653828772 $T=162340 150320 0 0 $X=160830 $Y=149290
X572 7 8 7 4 pe3_CDNS_724653828773 $T=138060 190125 0 0 $X=136550 $Y=189095
X573 8 2 7 4 pe3_CDNS_724653828773 $T=147620 190125 0 0 $X=146110 $Y=189095
X574 10 18 4 rpp1k1_3_CDNS_724653828774 $T=87870 117335 0 0 $X=82710 $Y=117115
X575 1 5 5 4 ne3_CDNS_724653828775 $T=17545 54415 0 0 $X=16745 $Y=54015
X576 3 5 6 4 ne3_CDNS_724653828775 $T=42480 54195 0 0 $X=41680 $Y=53795
X577 7 16 11 7 7 4 MASCO__A1 $T=216005 174905 0 0 $X=216005 $Y=174905
X578 7 16 12 7 7 4 MASCO__A1 $T=216005 194925 0 0 $X=216005 $Y=194925
X579 7 7 15 7 15 4 MASCO__A2 $T=10500 171290 0 0 $X=10500 $Y=171290
X580 7 7 16 7 15 4 MASCO__A2 $T=10500 188970 0 0 $X=10500 $Y=188970
X581 7 16 15 15 15 4 MASCO__A2 $T=32980 171290 0 0 $X=32980 $Y=171290
X582 7 15 16 15 15 4 MASCO__A2 $T=32980 188970 0 0 $X=32980 $Y=188970
X583 7 16 15 15 15 4 MASCO__A2 $T=55460 171290 0 0 $X=55460 $Y=171290
X584 7 15 16 15 15 4 MASCO__A2 $T=55460 188970 0 0 $X=55460 $Y=188970
X585 7 16 15 15 15 4 MASCO__A2 $T=77940 171290 0 0 $X=77940 $Y=171290
X586 7 15 16 15 15 4 MASCO__A2 $T=77940 188970 0 0 $X=77940 $Y=188970
X587 7 16 7 15 7 4 MASCO__A2 $T=100420 171290 0 0 $X=100420 $Y=171290
X588 7 15 7 15 7 4 MASCO__A2 $T=100420 188970 0 0 $X=100420 $Y=188970
X589 6 7 6 6 6 16 15 10 6 17
+ 4 MASCO__B5 $T=9330 114030 0 0 $X=9330 $Y=114030
X590 6 7 15 16 10 16 15 10 17 17
+ 4 MASCO__B5 $T=16130 114030 0 0 $X=16130 $Y=114030
X591 6 7 15 16 10 16 15 10 17 17
+ 4 MASCO__B5 $T=22930 114030 0 0 $X=22930 $Y=114030
X592 6 7 15 16 10 16 15 10 17 17
+ 4 MASCO__B5 $T=29730 114030 0 0 $X=29730 $Y=114030
X593 6 7 15 16 10 16 15 10 17 17
+ 4 MASCO__B5 $T=36530 114030 0 0 $X=36530 $Y=114030
X594 6 7 15 16 10 16 15 10 17 17
+ 4 MASCO__B5 $T=43330 114030 0 0 $X=43330 $Y=114030
X595 6 7 15 16 10 16 15 10 17 17
+ 4 MASCO__B5 $T=50130 114030 0 0 $X=50130 $Y=114030
X596 6 7 15 16 10 6 6 6 17 6
+ 4 MASCO__B5 $T=56930 114030 0 0 $X=56930 $Y=114030
X597 7 7 7 16 11 12 9 4 MASCO__A6 $T=164165 174905 0 0 $X=164165 $Y=174905
X598 7 7 7 16 12 9 11 4 MASCO__A6 $T=164165 194925 0 0 $X=164165 $Y=194925
X599 7 16 11 16 9 12 9 4 MASCO__A6 $T=177125 174905 0 0 $X=177125 $Y=174905
X600 7 16 12 16 12 9 11 4 MASCO__A6 $T=177125 194925 0 0 $X=177125 $Y=194925
X601 7 16 11 16 9 12 9 4 MASCO__A6 $T=190085 174905 0 0 $X=190085 $Y=174905
X602 7 16 9 16 12 9 11 4 MASCO__A6 $T=190085 194925 0 0 $X=190085 $Y=194925
X603 7 16 11 16 11 12 9 4 MASCO__A6 $T=203045 174905 0 0 $X=203045 $Y=174905
X604 7 16 9 16 12 9 11 4 MASCO__A6 $T=203045 194925 0 0 $X=203045 $Y=194925
X605 14 4 4 MOSVC3 w=3e-05 l=3e-05 $X=85530 $Y=8110 $dt=3
X606 14 4 4 MOSVC3 w=3e-05 l=3e-05 $X=85530 $Y=39350 $dt=3
X607 14 4 4 MOSVC3 w=3e-05 l=3e-05 $X=85530 $Y=70590 $dt=3
X608 13 4 4 MOSVC3 w=3e-05 l=3e-05 $X=122495 $Y=8050 $dt=3
X609 13 4 4 MOSVC3 w=3e-05 l=3e-05 $X=122495 $Y=39290 $dt=3
X610 13 4 4 MOSVC3 w=3e-05 l=3e-05 $X=122495 $Y=70530 $dt=3
D6 4 7 p_dnw AREA=2.36318e-09 PJ=0.00033402 perimeter=0.00033402 $X=4385 $Y=163650 $dt=4
D7 4 7 p_dnw AREA=2.57209e-10 PJ=8.388e-05 perimeter=8.388e-05 $X=134410 $Y=183535 $dt=4
D8 4 7 p_dnw AREA=1.81014e-09 PJ=0.00023539 perimeter=0.00023539 $X=158410 $Y=166295 $dt=4
D9 4 7 p_dnw AREA=8.15582e-10 PJ=0.0001871 perimeter=0.0001871 $X=158690 $Y=143730 $dt=4
D10 4 7 p_dnw AREA=9.45702e-09 PJ=0.00040696 perimeter=0.00040696 $X=159475 $Y=6005 $dt=4
D11 4 7 p_ddnw AREA=1.66704e-09 PJ=0.0001998 perimeter=0.0001998 $X=8060 $Y=112760 $dt=5
D12 6 7 p_dipdnwmv AREA=9.57098e-10 PJ=0.000169 perimeter=0.000169 $X=11910 $Y=116610 $dt=6
D13 4 7 p_dnw3 AREA=1.37701e-09 PJ=0 perimeter=0 $X=10500 $Y=171290 $dt=7
D14 4 7 p_dnw3 AREA=1.37701e-09 PJ=0 perimeter=0 $X=10500 $Y=188970 $dt=7
D15 4 4 p_dnw3 AREA=2.03309e-10 PJ=0.00024988 perimeter=0.00024988 $X=85100 $Y=7310 $dt=7
D16 4 4 p_dnw3 AREA=2.03309e-10 PJ=0.00024988 perimeter=0.00024988 $X=122065 $Y=7250 $dt=7
D17 4 7 p_dnw3 AREA=7.24806e-10 PJ=0 perimeter=0 $X=164165 $Y=174905 $dt=7
D18 4 7 p_dnw3 AREA=7.24806e-10 PJ=0 perimeter=0 $X=164165 $Y=194925 $dt=7
C19 16 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=161615 $Y=8145 $dt=9
C20 16 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=161615 $Y=39745 $dt=9
C21 16 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=161615 $Y=71345 $dt=9
C22 16 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=161615 $Y=102945 $dt=9
C23 16 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=196615 $Y=8145 $dt=9
C24 16 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=196615 $Y=39745 $dt=9
C25 16 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=196615 $Y=71345 $dt=9
C26 16 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=196615 $Y=102945 $dt=9
.ends ref_bias
