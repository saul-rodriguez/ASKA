************************************************************************
* auCdl Netlist:
* 
* Library Name:  CURRENT_SOURCE
* Top Cell Name: current_source_gm_10_en_r
* View Name:     schematic
* Netlisted on:  Aug 13 03:37:08 2024
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.LDD
*.SCALE METER
.PARAM



************************************************************************
* Library Name: CURRENT_SOURCE
* Cell Name:    current_source_gm_10_en_r
* View Name:    schematic
************************************************************************

.SUBCKT current_source_gm_10_en_r BIAS EN FB GNDA GNDHV IN OUT PACTIVE VDD3A 
+ VDDHV VSUBHV
*.PININFO BIAS:B EN:B FB:B GNDA:B GNDHV:B IN:B OUT:B PACTIVE:B VDD3A:B VDDHV:B 
*.PININFO VSUBHV:B
XC0 VDD3A GNDA GNDA / mosvc3 W=20u L=30u M=4.0 par1=4.0
MM30 VDD3A VDD3A VDD3A VDD3A PE3 W=10u L=5u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM26 net16 EN VDD3A VDD3A PE3 W=3u L=300n M=2.0 AD=2.88e-12 AS=2.88e-12 
+ PD=1.296e-05 PS=1.296e-05 NRD=0.045 NRS=0.045
MM35 net13 PACTIVE VDD3A VDD3A PE3 W=3u L=300n M=2.0 AD=2.88e-12 AS=2.88e-12 
+ PD=1.296e-05 PS=1.296e-05 NRD=0.045 NRS=0.045
MM23 net15 net15 VDD3A VDD3A PE3 W=10u L=1u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM29 VDD3A VDD3A VDD3A VDD3A PE3 W=10u L=5u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM11 net10 net4 VDD3A VDD3A PE3 W=10u L=5u M=2.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM9 net6 net4 VDD3A VDD3A PE3 W=10u L=5u M=2.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM10 net8 net4 VDD3A VDD3A PE3 W=10u L=5u M=20.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM20 VB net15 VDD3A VDD3A PE3 W=10u L=1u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM5 net9 net10 net8 VDD3A PE3 W=10u L=5u M=14.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM3 net7 net6 net8 VDD3A PE3 W=10u L=5u M=14.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM12 net4 net4 VDD3A VDD3A PE3 W=10u L=5u M=2.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM8 GNDA IN net6 net6 PE3 W=10u L=5u M=18.0 AD=2.93333e-12 AS=2.93333e-12 
+ PD=1.16978e-05 PS=1.16978e-05 NRD=0.027 NRS=0.027
MM7 GNDA net1 net10 net10 PE3 W=10u L=5u M=18.0 AD=2.93333e-12 AS=2.93333e-12 
+ PD=1.16978e-05 PS=1.16978e-05 NRD=0.027 NRS=0.027
MM25 net16 EN GNDA GNDA NE3 W=2u L=350.0n M=1.0 AD=9.6e-13 AS=9.6e-13 
+ PD=4.96e-06 PS=4.96e-06 NRD=0.135 NRS=0.135
MM24 net12 net16 GNDA GNDA NE3 W=5u L=350.0n M=4.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM34 net13 PACTIVE GNDA GNDA NE3 W=2u L=350.0n M=1.0 AD=9.6e-13 AS=9.6e-13 
+ PD=4.96e-06 PS=4.96e-06 NRD=0.135 NRS=0.135
MM32 net9 net13 GNDA GNDA NE3 W=5u L=350.0n M=4.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM22 net15 BIAS net14 GNDA NE3 W=10u L=10u M=2.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM21 net14 net12 GNDA GNDA NE3 W=10u L=10u M=2.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM19 net4 BIAS net5 GNDA NE3 W=10u L=10u M=2.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM18 BIAS BIAS net12 GNDA NE3 W=10u L=10u M=2.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM27 GNDA GNDA GNDA GNDA NE3 W=10u L=10u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM6 VB net9 GNDA GNDA NE3 W=5u L=500n M=4.0 AD=1.35e-12 AS=1.875e-12 
+ PD=5.54e-06 PS=8.25e-06 NRD=0.054 NRS=0.054
MM4 net7 net7 GNDA GNDA NE3 W=5u L=1u M=2.0 AD=2.4e-12 AS=2.4e-12 PD=1.096e-05 
+ PS=1.096e-05 NRD=0.054 NRS=0.054
MM2 net9 net7 GNDA GNDA NE3 W=5u L=1u M=2.0 AD=2.4e-12 AS=2.4e-12 PD=1.096e-05 
+ PS=1.096e-05 NRD=0.054 NRS=0.054
MM13 net5 net12 GNDA GNDA NE3 W=10u L=10u M=2.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM14 net12 net12 GNDA GNDA NE3 W=10u L=10u M=2.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM0 OUT VA FB VSUBHV NEDIA W=100.0000u L=1.25u M=8.0 $LDD[NEDIA]
MM1 VA VB GNDHV VSUBHV NEDIA W=50u L=1.25u M=1.0 $LDD[NEDIA]
RR1 VSUBHV GNDA 5.0 $[S_RES]
CC1 net9 net11 $[CMM5T] area=8.4e-10 perimeter=116.000000u M=7
RR7 GNDHV OUT 1.00618M $SUB=VSUBHV $[RPP1K1_3] $W=2u $L=2.04358m M=1
RR4 FB net1 5031.08 $SUB=GNDA $[RPP1K1_3] $W=2u $L=10u M=9
RR2 VA VDDHV 99.9954K $SUB=VSUBHV $[RPP1K1_3] $W=4u $L=411.22u M=1
RR3 GNDHV VA 25.0012K $SUB=VSUBHV $[RPP1K1_3] $W=4u $L=102.65u M=1
RR0 net11 VB 39.9966K $SUB=VDD3A $[RPP1K1_3] $W=4u $L=164.35u M=1
.ENDS


.SUBCKT mosvc3 G NW SB 
*.PININFO  G:B NW:B SB:B
.ENDS
