* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : dac6b_amp_n2                                 *
* Netlisted  : Wed Jun 26 14:49:12 2024                     *
* PVS Version: 23.10-p043 Mon Oct 2 18:09:08 PDT 2023      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(ne3) nem ndiff(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 1 MP(pe3) pem pdiff(D) p1trm(G) pdiff(S) nwtrm(B)
*.DEVTMPLT 2 NE3I_6() nemi_6 ndiff(D) p1trm(G) ndiff(S) pwitrm(B) dnwtrm(NW) bulk(SB)
*.DEVTMPLT 3 D(p_dnw) p_dnw bulk(POS) nwtrm(NEG)
*.DEVTMPLT 4 D(p_ddnw) p_ddnw bulk(POS) dnwtrm(NEG)
*.DEVTMPLT 5 D(p_dipdnwmv) p_dipwmv pwitrm(POS) dnwtrm(NEG)
*.DEVTMPLT 6 D(p_dnw3) p_dnwm bulk(POS) nwtrm(NEG)
*.DEVTMPLT 7 R(rpp1k1_3) rpp1k1_s p1trm(POS) p1trm(NEG) bulk(SUB)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_719427747080                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_719427747080 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_719427747080

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_719427747081                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_719427747081 1 2
** N=2 EP=2 FDC=0
.ends VIA1_C_CDNS_719427747081

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_719427747082                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_719427747082 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_719427747082

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_719427747083                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_719427747083 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_719427747083

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_719427747084                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_719427747084 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_719427747084

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_719427747085                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_719427747085 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_719427747085

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_719427747086                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_719427747086 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_719427747086

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_719427747087                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_719427747087 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_719427747087

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_719427747088                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_719427747088 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_719427747088

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_719427747089                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_719427747089 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_719427747089

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7194277470810                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7194277470810 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7194277470810

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7194277470811                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7194277470811 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7194277470811

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7194277470812                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7194277470812 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7194277470812

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7194277470813                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7194277470813 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7194277470813

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7194277470814                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7194277470814 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7194277470814

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7194277470816                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7194277470816 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7194277470816

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7194277470817                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7194277470817 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7194277470817

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7194277470818                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7194277470818 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7194277470818

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_7194277470819                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_7194277470819 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_7194277470819

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7194277470820                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7194277470820 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7194277470820

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7194277470822                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7194277470822 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7194277470822

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7194277470823                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7194277470823 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7194277470823

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7194277470824                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7194277470824 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7194277470824

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7194277470825                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7194277470825 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7194277470825

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7194277470826                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7194277470826 1 2
** N=2 EP=2 FDC=0
.ends VIA1_C_CDNS_7194277470826

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7194277470827                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7194277470827 1 2
** N=2 EP=2 FDC=0
.ends VIA2_C_CDNS_7194277470827

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7194277470828                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7194277470828 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7194277470828

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7194277470832                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7194277470832 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7194277470832

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7194277470833                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7194277470833 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7194277470833

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7194277470834                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7194277470834 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7194277470834

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_7194277470838                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_7194277470838 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_7194277470838

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_7194277470840                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_7194277470840 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_7194277470840

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_7194277470843                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_7194277470843 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_7194277470843

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7194277470846                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7194277470846 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7194277470846

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_719427747080                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_719427747080 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
M0 3 2 1 1 pe3 L=1e-05 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_719427747080

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_719427747081                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_719427747081 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
D1 5 4 p_dnw3 AREA=4.84812e-11 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=6
.ends pe3_CDNS_719427747081

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_719427747082                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_719427747082 1 2 3 4 5
** N=5 EP=5 FDC=3
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=1
D2 5 4 p_dnw3 AREA=6.70536e-11 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=6
.ends pe3_CDNS_719427747082

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_719427747083                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_719427747083 1 2 3 4 5
** N=5 EP=5 FDC=5
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=1
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=1
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=1
D4 5 4 p_dnw3 AREA=1.04198e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=6
.ends pe3_CDNS_719427747083

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_719427747084                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_719427747084 1 2 3 4 5
** N=5 EP=5 FDC=9
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=1
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=1
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=1
M4 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=6160 $Y=0 $dt=1
M5 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7700 $Y=0 $dt=1
M6 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=9240 $Y=0 $dt=1
M7 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=10780 $Y=0 $dt=1
D8 5 4 p_dnw3 AREA=1.78488e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=6
.ends pe3_CDNS_719427747084

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_719427747085                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_719427747085 1 2 3 4 5
** N=5 EP=5 FDC=17
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=1
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=1
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=1
M4 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=6160 $Y=0 $dt=1
M5 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7700 $Y=0 $dt=1
M6 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=9240 $Y=0 $dt=1
M7 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10780 $Y=0 $dt=1
M8 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12320 $Y=0 $dt=1
M9 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=13860 $Y=0 $dt=1
M10 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=15400 $Y=0 $dt=1
M11 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=16940 $Y=0 $dt=1
M12 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=18480 $Y=0 $dt=1
M13 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=20020 $Y=0 $dt=1
M14 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=21560 $Y=0 $dt=1
M15 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=23100 $Y=0 $dt=1
D16 5 4 p_dnw3 AREA=3.27067e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=6
.ends pe3_CDNS_719427747085

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_719427747086                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_719427747086 1 2 3 4 5
** N=5 EP=5 FDC=33
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=1
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=1
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=1
M4 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=6160 $Y=0 $dt=1
M5 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7700 $Y=0 $dt=1
M6 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=9240 $Y=0 $dt=1
M7 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10780 $Y=0 $dt=1
M8 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12320 $Y=0 $dt=1
M9 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=13860 $Y=0 $dt=1
M10 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=15400 $Y=0 $dt=1
M11 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=16940 $Y=0 $dt=1
M12 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=18480 $Y=0 $dt=1
M13 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=20020 $Y=0 $dt=1
M14 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=21560 $Y=0 $dt=1
M15 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=23100 $Y=0 $dt=1
M16 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=24640 $Y=0 $dt=1
M17 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=26180 $Y=0 $dt=1
M18 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=27720 $Y=0 $dt=1
M19 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=29260 $Y=0 $dt=1
M20 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=30800 $Y=0 $dt=1
M21 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=32340 $Y=0 $dt=1
M22 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=33880 $Y=0 $dt=1
M23 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=35420 $Y=0 $dt=1
M24 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=36960 $Y=0 $dt=1
M25 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=38500 $Y=0 $dt=1
M26 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=40040 $Y=0 $dt=1
M27 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=41580 $Y=0 $dt=1
M28 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=43120 $Y=0 $dt=1
M29 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=44660 $Y=0 $dt=1
M30 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=46200 $Y=0 $dt=1
M31 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=47740 $Y=0 $dt=1
D32 5 4 p_dnw3 AREA=6.24226e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=6
.ends pe3_CDNS_719427747086

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_719427747087                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_719427747087 1 2
** N=2 EP=2 FDC=1
R0 2 1 L=0.00021702 W=4e-06 $[rpp1k1_3] $SUB=2 $X=-4220 $Y=0 $dt=7
.ends rpp1k1_3_CDNS_719427747087

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_719427747088                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_719427747088 1 2 3 4 5
** N=5 EP=5 FDC=11
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=1
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=1
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=1
M4 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=6160 $Y=0 $dt=1
M5 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7700 $Y=0 $dt=1
M6 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=9240 $Y=0 $dt=1
M7 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10780 $Y=0 $dt=1
M8 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12320 $Y=0 $dt=1
M9 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=13860 $Y=0 $dt=1
D10 5 4 p_dnw3 AREA=2.15633e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=6
.ends pe3_CDNS_719427747088

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_719427747089                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_719427747089 1 2
** N=2 EP=2 FDC=1
R0 2 1 L=0.0008227 W=4e-06 $[rpp1k1_3] $SUB=2 $X=-4220 $Y=0 $dt=7
.ends rpp1k1_3_CDNS_719427747089

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7194277470810                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7194277470810 1 2 3
** N=3 EP=3 FDC=2
M0 2 2 1 1 pe3 L=2e-05 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
D1 3 1 p_dnw3 AREA=2.77621e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=6
.ends pe3_CDNS_7194277470810

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7194277470811                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7194277470811 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
M0 3 2 1 1 pe3 L=3e-07 W=6e-06 AD=2.88e-12 AS=2.88e-12 PD=1.296e-05 PS=1.296e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_7194277470811

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7194277470812                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7194277470812 1 2 3 4
** N=4 EP=4 FDC=3
M0 3 2 1 4 pe3 L=3.5e-07 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=3.5e-07 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=890 $Y=0 $dt=1
D2 3 4 p_dnw3 AREA=5.13756e-11 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=6
.ends pe3_CDNS_7194277470812

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7194277470813                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7194277470813 1 2 3 4
** N=4 EP=4 FDC=8
M0 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
M1 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=2540 $Y=0 $dt=0
M2 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=5080 $Y=0 $dt=0
M3 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7620 $Y=0 $dt=0
M4 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10160 $Y=0 $dt=0
M5 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12700 $Y=0 $dt=0
M6 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=15240 $Y=0 $dt=0
M7 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=17780 $Y=0 $dt=0
.ends ne3_CDNS_7194277470813

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7194277470815                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7194277470815 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=2e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
.ends ne3_CDNS_7194277470815

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7194277470816                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7194277470816 1 2
*.DEVICECLIMB
** N=2 EP=2 FDC=1
M0 1 1 1 1 pe3 L=1e-05 W=2e-06 AD=9.6e-13 AS=9.6e-13 PD=4.96e-06 PS=4.96e-06 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_7194277470816

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7194277470817                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7194277470817 1 2 3
** N=3 EP=3 FDC=4
M0 3 2 1 1 ne3 L=3.5e-07 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
M1 1 2 3 1 ne3 L=3.5e-07 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=890 $Y=0 $dt=0
M2 3 2 1 1 ne3 L=3.5e-07 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1780 $Y=0 $dt=0
M3 1 2 3 1 ne3 L=3.5e-07 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=2670 $Y=0 $dt=0
.ends ne3_CDNS_7194277470817

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7194277470818                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7194277470818 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=3.5e-07 W=2e-06 AD=9.6e-13 AS=9.6e-13 PD=4.96e-06 PS=4.96e-06 $X=0 $Y=0 $dt=0
.ends ne3_CDNS_7194277470818

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A1 1 2
*.DEVICECLIMB
** N=2 EP=2 FDC=2
X0 1 2 pe3_CDNS_7194277470816 $T=1510 3030 1 0 $X=0 $Y=0
X1 1 2 pe3_CDNS_7194277470816 $T=12750 3030 1 0 $X=11240 $Y=0
.ends MASCO__A1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A2 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 4 2 6 pe3_CDNS_719427747080 $T=1510 11030 1 0 $X=0 $Y=0
X1 1 5 3 6 pe3_CDNS_719427747080 $T=12750 11030 1 0 $X=11240 $Y=0
.ends MASCO__A2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3i_6_CDNS_7194277470814                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3i_6_CDNS_7194277470814 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=1
X0 1 2 3 1 4 5 NE3I_6 w=1e-05 l=2e-06 as=4.8e-12 ad=4.8e-12 ps=2.096e-05 pd=2.096e-05 $X=0 $Y=0 $dt=2
.ends ne3i_6_CDNS_7194277470814

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A3                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A3 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=2
X0 1 3 2 6 7 ne3i_6_CDNS_7194277470814 $T=4060 14570 1 0 $X=0 $Y=0
X1 1 5 4 6 7 ne3i_6_CDNS_7194277470814 $T=7460 14570 1 0 $X=3400 $Y=0
.ends MASCO__A3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A4                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A4 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=2
X0 1 5 4 6 7 ne3i_6_CDNS_7194277470814 $T=4060 4450 0 0 $X=0 $Y=0
X1 1 3 2 6 7 ne3i_6_CDNS_7194277470814 $T=7460 4450 0 0 $X=3400 $Y=0
.ends MASCO__A4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__B5                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__B5 1 2 3 4 5 6 7 8 9 10
+ 11
*.DEVICECLIMB
** N=11 EP=11 FDC=4
X0 1 3 10 5 9 2 11 MASCO__A3 $T=0 13180 0 0 $X=0 $Y=13180
X1 1 6 7 4 8 2 11 MASCO__A4 $T=0 0 0 0 $X=0 $Y=0
.ends MASCO__B5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A6                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A6 1 2 3 4 5 6 7 8
*.DEVICECLIMB
** N=8 EP=8 FDC=4
X0 1 2 4 7 3 8 MASCO__A2 $T=0 0 0 0 $X=0 $Y=0
X1 1 5 6 3 3 8 MASCO__A2 $T=22480 0 0 0 $X=22480 $Y=0
.ends MASCO__A6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: dac6b_amp_n2                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt dac6b_amp_n2 2 30 29 28 27 26 25 24 11 5
+ 22 23
** N=31 EP=12 FDC=372
X0 1 VIA1_C_CDNS_719427747080 $T=7445 56365 0 0 $X=7045 $Y=55655
X1 2 VIA1_C_CDNS_719427747080 $T=9985 58145 0 0 $X=9585 $Y=57435
X2 1 VIA1_C_CDNS_719427747080 $T=12525 56365 0 0 $X=12125 $Y=55655
X3 2 VIA1_C_CDNS_719427747080 $T=15065 58145 0 0 $X=14665 $Y=57435
X4 1 VIA1_C_CDNS_719427747080 $T=17605 56365 0 0 $X=17205 $Y=55655
X5 2 VIA1_C_CDNS_719427747080 $T=20145 58145 0 0 $X=19745 $Y=57435
X6 1 VIA1_C_CDNS_719427747080 $T=22685 56365 0 0 $X=22285 $Y=55655
X7 2 VIA1_C_CDNS_719427747080 $T=25225 58145 0 0 $X=24825 $Y=57435
X8 1 VIA1_C_CDNS_719427747080 $T=27765 56365 0 0 $X=27365 $Y=55655
X9 3 VIA1_C_CDNS_719427747080 $T=34200 58145 0 0 $X=33800 $Y=57435
X10 4 VIA1_C_CDNS_719427747080 $T=36740 56365 0 0 $X=36340 $Y=55655
X11 3 VIA1_C_CDNS_719427747080 $T=39280 58145 0 0 $X=38880 $Y=57435
X12 4 VIA1_C_CDNS_719427747080 $T=41820 56365 0 0 $X=41420 $Y=55655
X13 3 VIA1_C_CDNS_719427747080 $T=44360 58145 0 0 $X=43960 $Y=57435
X14 4 VIA1_C_CDNS_719427747080 $T=46900 56365 0 0 $X=46500 $Y=55655
X15 3 VIA1_C_CDNS_719427747080 $T=49440 58145 0 0 $X=49040 $Y=57435
X16 4 VIA1_C_CDNS_719427747080 $T=51980 56365 0 0 $X=51580 $Y=55655
X17 3 VIA1_C_CDNS_719427747080 $T=54520 58145 0 0 $X=54120 $Y=57435
X18 5 VIA1_C_CDNS_719427747080 $T=56070 146660 0 0 $X=55670 $Y=145950
X19 5 VIA1_C_CDNS_719427747080 $T=56070 173480 0 0 $X=55670 $Y=172770
X20 5 VIA1_C_CDNS_719427747080 $T=66380 146660 0 0 $X=65980 $Y=145950
X21 5 VIA1_C_CDNS_719427747080 $T=66380 173480 0 0 $X=65980 $Y=172770
X22 5 VIA1_C_CDNS_719427747080 $T=67540 146660 0 0 $X=67140 $Y=145950
X23 5 VIA1_C_CDNS_719427747080 $T=67540 173480 0 0 $X=67140 $Y=172770
X24 6 VIA1_C_CDNS_719427747080 $T=77620 144880 0 0 $X=77220 $Y=144170
X25 7 VIA1_C_CDNS_719427747080 $T=77620 175260 0 0 $X=77220 $Y=174550
X26 7 VIA1_C_CDNS_719427747080 $T=88860 143100 0 0 $X=88460 $Y=142390
X27 6 VIA1_C_CDNS_719427747080 $T=88860 177040 0 0 $X=88460 $Y=176330
X28 6 VIA1_C_CDNS_719427747080 $T=100100 144880 0 0 $X=99700 $Y=144170
X29 7 VIA1_C_CDNS_719427747080 $T=100100 175260 0 0 $X=99700 $Y=174550
X30 7 VIA1_C_CDNS_719427747080 $T=111340 143100 0 0 $X=110940 $Y=142390
X31 6 VIA1_C_CDNS_719427747080 $T=111340 177040 0 0 $X=110940 $Y=176330
X32 6 VIA1_C_CDNS_719427747080 $T=122580 144880 0 0 $X=122180 $Y=144170
X33 7 VIA1_C_CDNS_719427747080 $T=122580 175260 0 0 $X=122180 $Y=174550
X34 7 VIA1_C_CDNS_719427747080 $T=133820 143100 0 0 $X=133420 $Y=142390
X35 6 VIA1_C_CDNS_719427747080 $T=133820 177040 0 0 $X=133420 $Y=176330
X36 6 VIA1_C_CDNS_719427747080 $T=145060 144880 0 0 $X=144660 $Y=144170
X37 7 VIA1_C_CDNS_719427747080 $T=145060 175260 0 0 $X=144660 $Y=174550
X38 8 VIA1_C_CDNS_719427747080 $T=154405 72995 0 0 $X=154005 $Y=72285
X39 9 VIA1_C_CDNS_719427747080 $T=154405 94475 0 0 $X=154005 $Y=93765
X40 10 VIA1_C_CDNS_719427747080 $T=154405 115425 0 0 $X=154005 $Y=114715
X41 7 VIA1_C_CDNS_719427747080 $T=156300 143100 0 0 $X=155900 $Y=142390
X42 6 VIA1_C_CDNS_719427747080 $T=156300 177040 0 0 $X=155900 $Y=176330
X43 5 VIA1_C_CDNS_719427747080 $T=167770 146660 0 0 $X=167370 $Y=145950
X44 5 VIA1_C_CDNS_719427747080 $T=167770 173480 0 0 $X=167370 $Y=172770
X45 11 VIA1_C_CDNS_719427747080 $T=174945 74775 0 0 $X=174545 $Y=74065
X46 8 VIA1_C_CDNS_719427747080 $T=174945 96255 0 0 $X=174545 $Y=95545
X47 9 VIA1_C_CDNS_719427747080 $T=174945 117205 0 0 $X=174545 $Y=116495
X48 8 11 VIA1_C_CDNS_719427747081 $T=166585 72935 0 0 $X=155215 $Y=72795
X49 9 11 VIA1_C_CDNS_719427747081 $T=166585 94415 0 0 $X=155215 $Y=94275
X50 10 11 VIA1_C_CDNS_719427747081 $T=166585 115365 0 0 $X=155215 $Y=115225
X51 8 VIA1_C_CDNS_719427747082 $T=152520 72935 0 0 $X=151290 $Y=72795
X52 9 VIA1_C_CDNS_719427747082 $T=152520 94415 0 0 $X=151290 $Y=94275
X53 10 VIA1_C_CDNS_719427747082 $T=152520 115365 0 0 $X=151290 $Y=115225
X54 11 VIA1_C_CDNS_719427747083 $T=11260 15030 0 0 $X=11120 $Y=14320
X55 11 VIA1_C_CDNS_719427747083 $T=11260 39750 0 0 $X=11120 $Y=39040
X56 11 VIA1_C_CDNS_719427747083 $T=13800 15030 0 0 $X=13660 $Y=14320
X57 11 VIA1_C_CDNS_719427747083 $T=13800 39750 0 0 $X=13660 $Y=39040
X58 11 VIA1_C_CDNS_719427747083 $T=14500 15030 0 0 $X=14360 $Y=14320
X59 11 VIA1_C_CDNS_719427747083 $T=14500 39750 0 0 $X=14360 $Y=39040
X60 5 VIA1_C_CDNS_719427747083 $T=15440 146660 0 0 $X=15300 $Y=145950
X61 5 VIA1_C_CDNS_719427747083 $T=15440 173480 0 0 $X=15300 $Y=172770
X62 12 VIA1_C_CDNS_719427747083 $T=17040 11470 0 0 $X=16900 $Y=10760
X63 1 VIA1_C_CDNS_719427747083 $T=17040 41530 0 0 $X=16900 $Y=40820
X64 11 VIA1_C_CDNS_719427747083 $T=17740 15030 0 0 $X=17600 $Y=14320
X65 11 VIA1_C_CDNS_719427747083 $T=17740 39750 0 0 $X=17600 $Y=39040
X66 3 VIA1_C_CDNS_719427747083 $T=20280 13250 0 0 $X=20140 $Y=12540
X67 12 VIA1_C_CDNS_719427747083 $T=20280 43310 0 0 $X=20140 $Y=42600
X68 11 VIA1_C_CDNS_719427747083 $T=20980 15030 0 0 $X=20840 $Y=14320
X69 11 VIA1_C_CDNS_719427747083 $T=20980 39750 0 0 $X=20840 $Y=39040
X70 1 VIA1_C_CDNS_719427747083 $T=23520 9690 0 0 $X=23380 $Y=8980
X71 3 VIA1_C_CDNS_719427747083 $T=23520 45090 0 0 $X=23380 $Y=44380
X72 11 VIA1_C_CDNS_719427747083 $T=24220 15030 0 0 $X=24080 $Y=14320
X73 11 VIA1_C_CDNS_719427747083 $T=24220 39750 0 0 $X=24080 $Y=39040
X74 4 VIA1_C_CDNS_719427747083 $T=25980 144880 0 0 $X=25840 $Y=144170
X75 10 VIA1_C_CDNS_719427747083 $T=25980 175260 0 0 $X=25840 $Y=174550
X76 5 VIA1_C_CDNS_719427747083 $T=26680 146660 0 0 $X=26540 $Y=145950
X77 5 VIA1_C_CDNS_719427747083 $T=26680 173480 0 0 $X=26540 $Y=172770
X78 12 VIA1_C_CDNS_719427747083 $T=26760 11470 0 0 $X=26620 $Y=10760
X79 1 VIA1_C_CDNS_719427747083 $T=26760 41530 0 0 $X=26620 $Y=40820
X80 11 VIA1_C_CDNS_719427747083 $T=27460 15030 0 0 $X=27320 $Y=14320
X81 11 VIA1_C_CDNS_719427747083 $T=27460 39750 0 0 $X=27320 $Y=39040
X82 3 VIA1_C_CDNS_719427747083 $T=30000 13250 0 0 $X=29860 $Y=12540
X83 12 VIA1_C_CDNS_719427747083 $T=30000 43310 0 0 $X=29860 $Y=42600
X84 11 VIA1_C_CDNS_719427747083 $T=30700 15030 0 0 $X=30560 $Y=14320
X85 11 VIA1_C_CDNS_719427747083 $T=30700 39750 0 0 $X=30560 $Y=39040
X86 1 VIA1_C_CDNS_719427747083 $T=33240 9690 0 0 $X=33100 $Y=8980
X87 3 VIA1_C_CDNS_719427747083 $T=33240 45090 0 0 $X=33100 $Y=44380
X88 11 VIA1_C_CDNS_719427747083 $T=33940 15030 0 0 $X=33800 $Y=14320
X89 11 VIA1_C_CDNS_719427747083 $T=33940 39750 0 0 $X=33800 $Y=39040
X90 12 VIA1_C_CDNS_719427747083 $T=36480 11470 0 0 $X=36340 $Y=10760
X91 1 VIA1_C_CDNS_719427747083 $T=36480 41530 0 0 $X=36340 $Y=40820
X92 11 VIA1_C_CDNS_719427747083 $T=37180 15030 0 0 $X=37040 $Y=14320
X93 11 VIA1_C_CDNS_719427747083 $T=37180 39750 0 0 $X=37040 $Y=39040
X94 10 VIA1_C_CDNS_719427747083 $T=37220 143100 0 0 $X=37080 $Y=142390
X95 4 VIA1_C_CDNS_719427747083 $T=37220 177040 0 0 $X=37080 $Y=176330
X96 3 VIA1_C_CDNS_719427747083 $T=39720 13250 0 0 $X=39580 $Y=12540
X97 12 VIA1_C_CDNS_719427747083 $T=39720 43310 0 0 $X=39580 $Y=42600
X98 11 VIA1_C_CDNS_719427747083 $T=40420 15030 0 0 $X=40280 $Y=14320
X99 11 VIA1_C_CDNS_719427747083 $T=40420 39750 0 0 $X=40280 $Y=39040
X100 1 VIA1_C_CDNS_719427747083 $T=42960 9690 0 0 $X=42820 $Y=8980
X101 3 VIA1_C_CDNS_719427747083 $T=42960 45090 0 0 $X=42820 $Y=44380
X102 11 VIA1_C_CDNS_719427747083 $T=43660 15030 0 0 $X=43520 $Y=14320
X103 11 VIA1_C_CDNS_719427747083 $T=43660 39750 0 0 $X=43520 $Y=39040
X104 12 VIA1_C_CDNS_719427747083 $T=46200 11470 0 0 $X=46060 $Y=10760
X105 1 VIA1_C_CDNS_719427747083 $T=46200 41530 0 0 $X=46060 $Y=40820
X106 11 VIA1_C_CDNS_719427747083 $T=46900 15030 0 0 $X=46760 $Y=14320
X107 11 VIA1_C_CDNS_719427747083 $T=46900 39750 0 0 $X=46760 $Y=39040
X108 3 VIA1_C_CDNS_719427747083 $T=49440 13250 0 0 $X=49300 $Y=12540
X109 12 VIA1_C_CDNS_719427747083 $T=49440 43310 0 0 $X=49300 $Y=42600
X110 11 VIA1_C_CDNS_719427747083 $T=50140 15030 0 0 $X=50000 $Y=14320
X111 11 VIA1_C_CDNS_719427747083 $T=50140 39750 0 0 $X=50000 $Y=39040
X112 1 VIA1_C_CDNS_719427747083 $T=52680 9690 0 0 $X=52540 $Y=8980
X113 3 VIA1_C_CDNS_719427747083 $T=52680 45090 0 0 $X=52540 $Y=44380
X114 11 VIA1_C_CDNS_719427747083 $T=53380 15030 0 0 $X=53240 $Y=14320
X115 11 VIA1_C_CDNS_719427747083 $T=53380 39750 0 0 $X=53240 $Y=39040
X116 11 VIA1_C_CDNS_719427747083 $T=55920 15030 0 0 $X=55780 $Y=14320
X117 11 VIA1_C_CDNS_719427747083 $T=55920 39750 0 0 $X=55780 $Y=39040
X118 11 VIA1_C_CDNS_719427747084 $T=8940 15030 0 0 $X=7970 $Y=14370
X119 11 VIA1_C_CDNS_719427747084 $T=8940 39750 0 0 $X=7970 $Y=39090
X120 5 VIA1_C_CDNS_719427747084 $T=12920 146660 0 0 $X=11950 $Y=146000
X121 5 VIA1_C_CDNS_719427747084 $T=12920 173480 0 0 $X=11950 $Y=172820
X122 5 VIA1_C_CDNS_719427747084 $T=39740 146660 0 0 $X=38770 $Y=146000
X123 5 VIA1_C_CDNS_719427747084 $T=39740 173480 0 0 $X=38770 $Y=172820
X124 5 VIA1_C_CDNS_719427747084 $T=53550 146660 0 0 $X=52580 $Y=146000
X125 5 VIA1_C_CDNS_719427747084 $T=53550 173480 0 0 $X=52580 $Y=172820
X126 11 VIA1_C_CDNS_719427747084 $T=57730 15030 0 0 $X=56760 $Y=14370
X127 11 VIA1_C_CDNS_719427747084 $T=57730 39750 0 0 $X=56760 $Y=39090
X128 5 VIA1_C_CDNS_719427747084 $T=170290 146660 0 0 $X=169320 $Y=146000
X129 5 VIA1_C_CDNS_719427747084 $T=170290 173480 0 0 $X=169320 $Y=172820
X130 11 VIA1_C_CDNS_719427747085 $T=10335 15030 0 0 $X=10195 $Y=14280
X131 11 VIA1_C_CDNS_719427747085 $T=10335 39750 0 0 $X=10195 $Y=39000
X132 2 VIA1_C_CDNS_719427747086 $T=8715 70535 0 0 $X=8315 $Y=70345
X133 2 VIA1_C_CDNS_719427747086 $T=11255 70535 0 0 $X=10855 $Y=70345
X134 2 VIA1_C_CDNS_719427747086 $T=13795 70535 0 0 $X=13395 $Y=70345
X135 1 VIA1_C_CDNS_719427747086 $T=15770 27420 0 0 $X=15370 $Y=27230
X136 2 VIA1_C_CDNS_719427747086 $T=16335 70535 0 0 $X=15935 $Y=70345
X137 2 VIA1_C_CDNS_719427747086 $T=18875 70535 0 0 $X=18475 $Y=70345
X138 1 VIA1_C_CDNS_719427747086 $T=19010 27420 0 0 $X=18610 $Y=27230
X139 4 VIA1_C_CDNS_719427747086 $T=20710 160140 0 0 $X=20310 $Y=159950
X140 2 VIA1_C_CDNS_719427747086 $T=21415 70535 0 0 $X=21015 $Y=70345
X141 1 VIA1_C_CDNS_719427747086 $T=22250 27420 0 0 $X=21850 $Y=27230
X142 2 VIA1_C_CDNS_719427747086 $T=23955 70535 0 0 $X=23555 $Y=70345
X143 1 VIA1_C_CDNS_719427747086 $T=25490 27420 0 0 $X=25090 $Y=27230
X144 2 VIA1_C_CDNS_719427747086 $T=26495 70535 0 0 $X=26095 $Y=70345
X145 1 VIA1_C_CDNS_719427747086 $T=28730 27420 0 0 $X=28330 $Y=27230
X146 4 VIA1_C_CDNS_719427747086 $T=31950 160140 0 0 $X=31550 $Y=159950
X147 1 VIA1_C_CDNS_719427747086 $T=31970 27420 0 0 $X=31570 $Y=27230
X148 1 VIA1_C_CDNS_719427747086 $T=35210 27420 0 0 $X=34810 $Y=27230
X149 2 VIA1_C_CDNS_719427747086 $T=35470 70535 0 0 $X=35070 $Y=70345
X150 2 VIA1_C_CDNS_719427747086 $T=38010 70535 0 0 $X=37610 $Y=70345
X151 1 VIA1_C_CDNS_719427747086 $T=38450 27420 0 0 $X=38050 $Y=27230
X152 2 VIA1_C_CDNS_719427747086 $T=40550 70535 0 0 $X=40150 $Y=70345
X153 1 VIA1_C_CDNS_719427747086 $T=41690 27420 0 0 $X=41290 $Y=27230
X154 2 VIA1_C_CDNS_719427747086 $T=43090 70535 0 0 $X=42690 $Y=70345
X155 1 VIA1_C_CDNS_719427747086 $T=44930 27420 0 0 $X=44530 $Y=27230
X156 2 VIA1_C_CDNS_719427747086 $T=45630 70535 0 0 $X=45230 $Y=70345
X157 1 VIA1_C_CDNS_719427747086 $T=48170 27420 0 0 $X=47770 $Y=27230
X158 2 VIA1_C_CDNS_719427747086 $T=48170 70535 0 0 $X=47770 $Y=70345
X159 2 VIA1_C_CDNS_719427747086 $T=50710 70535 0 0 $X=50310 $Y=70345
X160 1 VIA1_C_CDNS_719427747086 $T=51410 27420 0 0 $X=51010 $Y=27230
X161 2 VIA1_C_CDNS_719427747086 $T=53250 70535 0 0 $X=52850 $Y=70345
X162 2 VIA1_C_CDNS_719427747086 $T=63205 70535 0 0 $X=62805 $Y=70345
X163 2 VIA1_C_CDNS_719427747086 $T=65745 70535 0 0 $X=65345 $Y=70345
X164 2 VIA1_C_CDNS_719427747086 $T=68285 70535 0 0 $X=67885 $Y=70345
X165 2 VIA1_C_CDNS_719427747086 $T=70825 70535 0 0 $X=70425 $Y=70345
X166 6 VIA1_C_CDNS_719427747086 $T=72580 160140 0 0 $X=72180 $Y=159950
X167 2 VIA1_C_CDNS_719427747086 $T=73365 70535 0 0 $X=72965 $Y=70345
X168 2 VIA1_C_CDNS_719427747086 $T=75905 70535 0 0 $X=75505 $Y=70345
X169 2 VIA1_C_CDNS_719427747086 $T=78445 70535 0 0 $X=78045 $Y=70345
X170 2 VIA1_C_CDNS_719427747086 $T=80985 70535 0 0 $X=80585 $Y=70345
X171 6 VIA1_C_CDNS_719427747086 $T=83820 160140 0 0 $X=83420 $Y=159950
X172 6 VIA1_C_CDNS_719427747086 $T=95060 160140 0 0 $X=94660 $Y=159950
X173 6 VIA1_C_CDNS_719427747086 $T=106300 160140 0 0 $X=105900 $Y=159950
X174 6 VIA1_C_CDNS_719427747086 $T=117540 160140 0 0 $X=117140 $Y=159950
X175 6 VIA1_C_CDNS_719427747086 $T=128780 160140 0 0 $X=128380 $Y=159950
X176 6 VIA1_C_CDNS_719427747086 $T=140020 160140 0 0 $X=139620 $Y=159950
X177 6 VIA1_C_CDNS_719427747086 $T=151260 160140 0 0 $X=150860 $Y=159950
X178 9 VIA1_C_CDNS_719427747086 $T=224435 24760 1 0 $X=224035 $Y=24570
X179 9 VIA1_C_CDNS_719427747086 $T=225975 24760 1 0 $X=225575 $Y=24570
X180 9 VIA1_C_CDNS_719427747086 $T=227515 24760 1 0 $X=227115 $Y=24570
X181 9 VIA1_C_CDNS_719427747086 $T=229055 24760 1 0 $X=228655 $Y=24570
X182 9 VIA1_C_CDNS_719427747086 $T=230595 24760 1 0 $X=230195 $Y=24570
X183 9 VIA1_C_CDNS_719427747086 $T=232135 24760 1 0 $X=231735 $Y=24570
X184 9 VIA1_C_CDNS_719427747086 $T=233675 24760 1 0 $X=233275 $Y=24570
X185 9 VIA1_C_CDNS_719427747086 $T=235215 24760 1 0 $X=234815 $Y=24570
X186 9 VIA1_C_CDNS_719427747086 $T=236755 24760 1 0 $X=236355 $Y=24570
X187 9 VIA1_C_CDNS_719427747086 $T=238295 24760 1 0 $X=237895 $Y=24570
X188 9 VIA1_C_CDNS_719427747086 $T=247255 24760 1 0 $X=246855 $Y=24570
X189 9 VIA1_C_CDNS_719427747086 $T=248795 24760 1 0 $X=248395 $Y=24570
X190 9 VIA1_C_CDNS_719427747086 $T=250335 24760 1 0 $X=249935 $Y=24570
X191 9 VIA1_C_CDNS_719427747086 $T=251875 24760 1 0 $X=251475 $Y=24570
X192 9 VIA1_C_CDNS_719427747086 $T=253415 24760 1 0 $X=253015 $Y=24570
X193 9 VIA1_C_CDNS_719427747086 $T=254955 24760 1 0 $X=254555 $Y=24570
X194 9 VIA1_C_CDNS_719427747086 $T=256495 24760 1 0 $X=256095 $Y=24570
X195 9 VIA1_C_CDNS_719427747086 $T=258035 24760 1 0 $X=257635 $Y=24570
X196 9 VIA1_C_CDNS_719427747086 $T=259575 24760 1 0 $X=259175 $Y=24570
X197 9 VIA1_C_CDNS_719427747086 $T=261115 24760 1 0 $X=260715 $Y=24570
X198 9 VIA1_C_CDNS_719427747086 $T=262655 24760 1 0 $X=262255 $Y=24570
X199 9 VIA1_C_CDNS_719427747086 $T=264195 24760 1 0 $X=263795 $Y=24570
X200 9 VIA1_C_CDNS_719427747086 $T=265735 24760 1 0 $X=265335 $Y=24570
X201 9 VIA1_C_CDNS_719427747086 $T=267275 24760 1 0 $X=266875 $Y=24570
X202 9 VIA1_C_CDNS_719427747086 $T=268815 24760 1 0 $X=268415 $Y=24570
X203 9 VIA1_C_CDNS_719427747086 $T=270355 24760 1 0 $X=269955 $Y=24570
X204 9 VIA1_C_CDNS_719427747086 $T=271895 24760 1 0 $X=271495 $Y=24570
X205 9 VIA1_C_CDNS_719427747086 $T=273435 24760 1 0 $X=273035 $Y=24570
X206 9 VIA1_C_CDNS_719427747086 $T=274975 24760 1 0 $X=274575 $Y=24570
X207 9 VIA1_C_CDNS_719427747086 $T=276515 24760 1 0 $X=276115 $Y=24570
X208 9 VIA1_C_CDNS_719427747086 $T=278055 24760 1 0 $X=277655 $Y=24570
X209 9 VIA1_C_CDNS_719427747086 $T=279595 24760 1 0 $X=279195 $Y=24570
X210 9 VIA1_C_CDNS_719427747086 $T=281135 24760 1 0 $X=280735 $Y=24570
X211 9 VIA1_C_CDNS_719427747086 $T=282675 24760 1 0 $X=282275 $Y=24570
X212 9 VIA1_C_CDNS_719427747086 $T=284215 24760 1 0 $X=283815 $Y=24570
X213 9 VIA1_C_CDNS_719427747086 $T=285755 24760 1 0 $X=285355 $Y=24570
X214 9 VIA1_C_CDNS_719427747086 $T=287295 24760 1 0 $X=286895 $Y=24570
X215 9 VIA1_C_CDNS_719427747086 $T=288835 24760 1 0 $X=288435 $Y=24570
X216 9 VIA1_C_CDNS_719427747086 $T=290375 24760 1 0 $X=289975 $Y=24570
X217 9 VIA1_C_CDNS_719427747086 $T=291915 24760 1 0 $X=291515 $Y=24570
X218 9 VIA1_C_CDNS_719427747086 $T=293455 24760 1 0 $X=293055 $Y=24570
X219 9 VIA1_C_CDNS_719427747086 $T=294995 24760 1 0 $X=294595 $Y=24570
X220 9 VIA1_C_CDNS_719427747086 $T=303070 24760 1 0 $X=302670 $Y=24570
X221 9 VIA1_C_CDNS_719427747086 $T=304610 24760 1 0 $X=304210 $Y=24570
X222 9 VIA1_C_CDNS_719427747086 $T=306150 24760 1 0 $X=305750 $Y=24570
X223 9 VIA1_C_CDNS_719427747086 $T=307690 24760 1 0 $X=307290 $Y=24570
X224 9 VIA1_C_CDNS_719427747086 $T=309230 24760 1 0 $X=308830 $Y=24570
X225 9 VIA1_C_CDNS_719427747086 $T=310770 24760 1 0 $X=310370 $Y=24570
X226 9 VIA1_C_CDNS_719427747086 $T=312310 24760 1 0 $X=311910 $Y=24570
X227 9 VIA1_C_CDNS_719427747086 $T=313850 24760 1 0 $X=313450 $Y=24570
X228 9 VIA1_C_CDNS_719427747086 $T=315390 24760 1 0 $X=314990 $Y=24570
X229 9 VIA1_C_CDNS_719427747086 $T=316930 24760 1 0 $X=316530 $Y=24570
X230 9 VIA1_C_CDNS_719427747086 $T=318470 24760 1 0 $X=318070 $Y=24570
X231 9 VIA1_C_CDNS_719427747086 $T=320010 24760 1 0 $X=319610 $Y=24570
X232 9 VIA1_C_CDNS_719427747086 $T=321550 24760 1 0 $X=321150 $Y=24570
X233 9 VIA1_C_CDNS_719427747086 $T=323090 24760 1 0 $X=322690 $Y=24570
X234 9 VIA1_C_CDNS_719427747086 $T=324630 24760 1 0 $X=324230 $Y=24570
X235 9 VIA1_C_CDNS_719427747086 $T=326170 24760 1 0 $X=325770 $Y=24570
X236 9 VIA1_C_CDNS_719427747086 $T=333835 24760 1 0 $X=333435 $Y=24570
X237 9 VIA1_C_CDNS_719427747086 $T=335375 24760 1 0 $X=334975 $Y=24570
X238 9 VIA1_C_CDNS_719427747086 $T=336915 24760 1 0 $X=336515 $Y=24570
X239 9 VIA1_C_CDNS_719427747086 $T=338455 24760 1 0 $X=338055 $Y=24570
X240 9 VIA1_C_CDNS_719427747086 $T=339995 24760 1 0 $X=339595 $Y=24570
X241 9 VIA1_C_CDNS_719427747086 $T=341535 24760 1 0 $X=341135 $Y=24570
X242 9 VIA1_C_CDNS_719427747086 $T=343075 24760 1 0 $X=342675 $Y=24570
X243 9 VIA1_C_CDNS_719427747086 $T=344615 24760 1 0 $X=344215 $Y=24570
X244 9 VIA1_C_CDNS_719427747086 $T=352300 24760 1 0 $X=351900 $Y=24570
X245 9 VIA1_C_CDNS_719427747086 $T=353840 24760 1 0 $X=353440 $Y=24570
X246 9 VIA1_C_CDNS_719427747086 $T=355380 24760 1 0 $X=354980 $Y=24570
X247 9 VIA1_C_CDNS_719427747086 $T=356920 24760 1 0 $X=356520 $Y=24570
X248 9 VIA1_C_CDNS_719427747086 $T=364635 24760 1 0 $X=364235 $Y=24570
X249 9 VIA1_C_CDNS_719427747086 $T=366175 24760 1 0 $X=365775 $Y=24570
X250 9 VIA1_C_CDNS_719427747086 $T=374010 24760 1 0 $X=373610 $Y=24570
X251 1 VIA2_C_CDNS_719427747087 $T=6660 9690 0 0 $X=5690 $Y=9030
X252 1 VIA2_C_CDNS_719427747087 $T=6660 41530 0 0 $X=5690 $Y=40870
X253 6 VIA2_C_CDNS_719427747087 $T=51270 144880 0 0 $X=50300 $Y=144220
X254 6 VIA2_C_CDNS_719427747087 $T=51270 177040 0 0 $X=50300 $Y=176380
X255 3 VIA2_C_CDNS_719427747087 $T=60010 13250 0 0 $X=59040 $Y=12590
X256 3 VIA2_C_CDNS_719427747087 $T=60010 45090 0 0 $X=59040 $Y=44430
X257 12 VIA2_C_CDNS_719427747087 $T=62290 11470 0 0 $X=61320 $Y=10810
X258 12 VIA2_C_CDNS_719427747087 $T=62290 43310 0 0 $X=61320 $Y=42650
X259 7 VIA2_C_CDNS_719427747087 $T=172570 143100 0 0 $X=171600 $Y=142440
X260 7 VIA2_C_CDNS_719427747087 $T=172570 175260 0 0 $X=171600 $Y=174600
X261 1 VIA2_C_CDNS_719427747088 $T=6660 27420 0 0 $X=5690 $Y=27280
X262 6 VIA2_C_CDNS_719427747088 $T=51270 160140 0 0 $X=50300 $Y=160000
X263 12 VIA1_C_CDNS_719427747089 $T=61935 55475 0 0 $X=61795 $Y=54505
X264 13 VIA1_C_CDNS_719427747089 $T=64475 57755 0 0 $X=64335 $Y=56785
X265 12 VIA1_C_CDNS_719427747089 $T=67015 55475 0 0 $X=66875 $Y=54505
X266 13 VIA1_C_CDNS_719427747089 $T=69555 57755 0 0 $X=69415 $Y=56785
X267 12 VIA1_C_CDNS_719427747089 $T=72095 55475 0 0 $X=71955 $Y=54505
X268 13 VIA1_C_CDNS_719427747089 $T=74635 57755 0 0 $X=74495 $Y=56785
X269 12 VIA1_C_CDNS_719427747089 $T=77175 55475 0 0 $X=77035 $Y=54505
X270 13 VIA1_C_CDNS_719427747089 $T=79715 57755 0 0 $X=79575 $Y=56785
X271 12 VIA1_C_CDNS_719427747089 $T=82255 55475 0 0 $X=82115 $Y=54505
X272 5 VIA1_C_CDNS_7194277470810 $T=214955 116235 0 0 $X=213985 $Y=116095
X273 5 VIA1_C_CDNS_7194277470810 $T=217155 78635 0 0 $X=216185 $Y=78495
X274 5 VIA1_C_CDNS_7194277470810 $T=217155 97435 0 0 $X=216185 $Y=97295
X275 5 VIA1_C_CDNS_7194277470810 $T=217155 116235 0 0 $X=216185 $Y=116095
X276 5 VIA1_C_CDNS_7194277470810 $T=217155 135035 0 0 $X=216185 $Y=134895
X277 5 VIA1_C_CDNS_7194277470810 $T=217155 153835 0 0 $X=216185 $Y=153695
X278 14 VIA1_C_CDNS_7194277470810 $T=226195 114675 0 0 $X=225225 $Y=114535
X279 5 VIA1_C_CDNS_7194277470810 $T=229015 78635 0 0 $X=228045 $Y=78495
X280 5 VIA1_C_CDNS_7194277470810 $T=229015 97435 0 0 $X=228045 $Y=97295
X281 5 VIA1_C_CDNS_7194277470810 $T=229015 116235 0 0 $X=228045 $Y=116095
X282 5 VIA1_C_CDNS_7194277470810 $T=229015 135035 0 0 $X=228045 $Y=134895
X283 5 VIA1_C_CDNS_7194277470810 $T=229015 153835 0 0 $X=228045 $Y=153695
X284 15 VIA1_C_CDNS_7194277470810 $T=237385 113895 0 0 $X=236415 $Y=113755
X285 5 VIA1_C_CDNS_7194277470810 $T=240255 78635 0 0 $X=239285 $Y=78495
X286 5 VIA1_C_CDNS_7194277470810 $T=240255 97435 0 0 $X=239285 $Y=97295
X287 5 VIA1_C_CDNS_7194277470810 $T=240255 116235 0 0 $X=239285 $Y=116095
X288 5 VIA1_C_CDNS_7194277470810 $T=240255 135035 0 0 $X=239285 $Y=134895
X289 5 VIA1_C_CDNS_7194277470810 $T=240255 153835 0 0 $X=239285 $Y=153695
X290 16 VIA1_C_CDNS_7194277470810 $T=248625 113115 0 0 $X=247655 $Y=112975
X291 5 VIA1_C_CDNS_7194277470810 $T=251495 78635 0 0 $X=250525 $Y=78495
X292 5 VIA1_C_CDNS_7194277470810 $T=251495 97435 0 0 $X=250525 $Y=97295
X293 5 VIA1_C_CDNS_7194277470810 $T=251495 116235 0 0 $X=250525 $Y=116095
X294 5 VIA1_C_CDNS_7194277470810 $T=251495 135035 0 0 $X=250525 $Y=134895
X295 5 VIA1_C_CDNS_7194277470810 $T=251495 153835 0 0 $X=250525 $Y=153695
X296 17 VIA1_C_CDNS_7194277470810 $T=259865 111555 0 0 $X=258895 $Y=111415
X297 5 VIA1_C_CDNS_7194277470810 $T=262735 78635 0 0 $X=261765 $Y=78495
X298 5 VIA1_C_CDNS_7194277470810 $T=262735 97435 0 0 $X=261765 $Y=97295
X299 5 VIA1_C_CDNS_7194277470810 $T=262735 116235 0 0 $X=261765 $Y=116095
X300 5 VIA1_C_CDNS_7194277470810 $T=262735 135035 0 0 $X=261765 $Y=134895
X301 5 VIA1_C_CDNS_7194277470810 $T=262735 153835 0 0 $X=261765 $Y=153695
X302 18 VIA1_C_CDNS_7194277470810 $T=271105 115455 0 0 $X=270135 $Y=115315
X303 5 VIA1_C_CDNS_7194277470810 $T=273975 78635 0 0 $X=273005 $Y=78495
X304 5 VIA1_C_CDNS_7194277470810 $T=273975 97435 0 0 $X=273005 $Y=97295
X305 5 VIA1_C_CDNS_7194277470810 $T=273975 116235 0 0 $X=273005 $Y=116095
X306 5 VIA1_C_CDNS_7194277470810 $T=273975 135035 0 0 $X=273005 $Y=134895
X307 5 VIA1_C_CDNS_7194277470810 $T=273975 153835 0 0 $X=273005 $Y=153695
X308 19 VIA1_C_CDNS_7194277470810 $T=282345 109995 0 0 $X=281375 $Y=109855
X309 5 VIA1_C_CDNS_7194277470810 $T=285215 78635 0 0 $X=284245 $Y=78495
X310 5 VIA1_C_CDNS_7194277470810 $T=285215 97435 0 0 $X=284245 $Y=97295
X311 5 VIA1_C_CDNS_7194277470810 $T=285215 116235 0 0 $X=284245 $Y=116095
X312 5 VIA1_C_CDNS_7194277470810 $T=285215 135035 0 0 $X=284245 $Y=134895
X313 5 VIA1_C_CDNS_7194277470810 $T=285215 153835 0 0 $X=284245 $Y=153695
X314 18 VIA1_C_CDNS_7194277470810 $T=293585 115455 0 0 $X=292615 $Y=115315
X315 5 VIA1_C_CDNS_7194277470810 $T=296455 78635 0 0 $X=295485 $Y=78495
X316 5 VIA1_C_CDNS_7194277470810 $T=296455 97435 0 0 $X=295485 $Y=97295
X317 5 VIA1_C_CDNS_7194277470810 $T=296455 116235 0 0 $X=295485 $Y=116095
X318 5 VIA1_C_CDNS_7194277470810 $T=296455 135035 0 0 $X=295485 $Y=134895
X319 5 VIA1_C_CDNS_7194277470810 $T=296455 153835 0 0 $X=295485 $Y=153695
X320 16 VIA1_C_CDNS_7194277470810 $T=304825 113115 0 0 $X=303855 $Y=112975
X321 5 VIA1_C_CDNS_7194277470810 $T=307695 78635 0 0 $X=306725 $Y=78495
X322 5 VIA1_C_CDNS_7194277470810 $T=307695 97435 0 0 $X=306725 $Y=97295
X323 5 VIA1_C_CDNS_7194277470810 $T=307695 116235 0 0 $X=306725 $Y=116095
X324 5 VIA1_C_CDNS_7194277470810 $T=307695 135035 0 0 $X=306725 $Y=134895
X325 5 VIA1_C_CDNS_7194277470810 $T=307695 153835 0 0 $X=306725 $Y=153695
X326 15 VIA1_C_CDNS_7194277470810 $T=316065 113895 0 0 $X=315095 $Y=113755
X327 5 VIA1_C_CDNS_7194277470810 $T=318315 78635 0 0 $X=317345 $Y=78495
X328 5 VIA1_C_CDNS_7194277470810 $T=318935 97435 0 0 $X=317965 $Y=97295
X329 5 VIA1_C_CDNS_7194277470810 $T=318935 116235 0 0 $X=317965 $Y=116095
X330 5 VIA1_C_CDNS_7194277470810 $T=318935 135035 0 0 $X=317965 $Y=134895
X331 5 VIA1_C_CDNS_7194277470810 $T=318935 153835 0 0 $X=317965 $Y=153695
X332 14 VIA1_C_CDNS_7194277470810 $T=327305 114675 0 0 $X=326335 $Y=114535
X333 5 VIA1_C_CDNS_7194277470810 $T=329555 78635 0 0 $X=328585 $Y=78495
X334 5 VIA1_C_CDNS_7194277470810 $T=330175 97435 0 0 $X=329205 $Y=97295
X335 5 VIA1_C_CDNS_7194277470810 $T=330175 116235 0 0 $X=329205 $Y=116095
X336 5 VIA1_C_CDNS_7194277470810 $T=330175 135035 0 0 $X=329205 $Y=134895
X337 5 VIA1_C_CDNS_7194277470810 $T=330175 153835 0 0 $X=329205 $Y=153695
X338 14 VIA1_C_CDNS_7194277470810 $T=338545 114675 0 0 $X=337575 $Y=114535
X339 5 VIA1_C_CDNS_7194277470810 $T=340795 78635 0 0 $X=339825 $Y=78495
X340 5 VIA1_C_CDNS_7194277470810 $T=341415 97435 0 0 $X=340445 $Y=97295
X341 5 VIA1_C_CDNS_7194277470810 $T=341415 116235 0 0 $X=340445 $Y=116095
X342 5 VIA1_C_CDNS_7194277470810 $T=341415 135035 0 0 $X=340445 $Y=134895
X343 5 VIA1_C_CDNS_7194277470810 $T=341415 153835 0 0 $X=340445 $Y=153695
X344 14 VIA1_C_CDNS_7194277470810 $T=349785 114675 0 0 $X=348815 $Y=114535
X345 5 VIA1_C_CDNS_7194277470810 $T=352035 78635 0 0 $X=351065 $Y=78495
X346 5 VIA1_C_CDNS_7194277470810 $T=352655 97435 0 0 $X=351685 $Y=97295
X347 5 VIA1_C_CDNS_7194277470810 $T=352655 116235 0 0 $X=351685 $Y=116095
X348 5 VIA1_C_CDNS_7194277470810 $T=352655 135035 0 0 $X=351685 $Y=134895
X349 5 VIA1_C_CDNS_7194277470810 $T=352655 153835 0 0 $X=351685 $Y=153695
X350 14 VIA1_C_CDNS_7194277470810 $T=361025 114675 0 0 $X=360055 $Y=114535
X351 5 VIA1_C_CDNS_7194277470810 $T=363275 78635 0 0 $X=362305 $Y=78495
X352 5 VIA1_C_CDNS_7194277470810 $T=363845 97435 0 0 $X=362875 $Y=97295
X353 5 VIA1_C_CDNS_7194277470810 $T=363845 116235 0 0 $X=362875 $Y=116095
X354 5 VIA1_C_CDNS_7194277470810 $T=363845 135035 0 0 $X=362875 $Y=134895
X355 5 VIA1_C_CDNS_7194277470810 $T=363845 153835 0 0 $X=362875 $Y=153695
X356 5 VIA1_C_CDNS_7194277470811 $T=205165 59835 0 0 $X=204245 $Y=59645
X357 5 VIA1_C_CDNS_7194277470811 $T=205165 78635 0 0 $X=204245 $Y=78445
X358 5 VIA1_C_CDNS_7194277470811 $T=205165 97435 0 0 $X=204245 $Y=97245
X359 5 VIA1_C_CDNS_7194277470811 $T=205165 116235 0 0 $X=204245 $Y=116045
X360 5 VIA1_C_CDNS_7194277470811 $T=205165 135035 0 0 $X=204245 $Y=134845
X361 5 VIA1_C_CDNS_7194277470811 $T=205165 153835 0 0 $X=204245 $Y=153645
X362 5 VIA1_C_CDNS_7194277470811 $T=205165 172635 0 0 $X=204245 $Y=172445
X363 5 VIA1_C_CDNS_7194277470811 $T=205165 177475 0 0 $X=204245 $Y=177285
X364 5 VIA1_C_CDNS_7194277470811 $T=210435 48755 0 0 $X=209515 $Y=48565
X365 5 VIA1_C_CDNS_7194277470811 $T=210435 59835 0 0 $X=209515 $Y=59645
X366 5 VIA1_C_CDNS_7194277470811 $T=210435 78635 0 0 $X=209515 $Y=78445
X367 5 VIA1_C_CDNS_7194277470811 $T=210435 97435 0 0 $X=209515 $Y=97245
X368 5 VIA1_C_CDNS_7194277470811 $T=210435 116235 0 0 $X=209515 $Y=116045
X369 5 VIA1_C_CDNS_7194277470811 $T=210435 135035 0 0 $X=209515 $Y=134845
X370 5 VIA1_C_CDNS_7194277470811 $T=210435 153835 0 0 $X=209515 $Y=153645
X371 5 VIA1_C_CDNS_7194277470811 $T=210435 172635 0 0 $X=209515 $Y=172445
X372 5 VIA1_C_CDNS_7194277470811 $T=214955 59835 0 0 $X=214035 $Y=59645
X373 5 VIA1_C_CDNS_7194277470811 $T=214955 78635 0 0 $X=214035 $Y=78445
X374 5 VIA1_C_CDNS_7194277470811 $T=214955 97435 0 0 $X=214035 $Y=97245
X375 5 VIA1_C_CDNS_7194277470811 $T=214955 135035 0 0 $X=214035 $Y=134845
X376 5 VIA1_C_CDNS_7194277470811 $T=214955 153835 0 0 $X=214035 $Y=153645
X377 5 VIA1_C_CDNS_7194277470811 $T=214955 172635 0 0 $X=214035 $Y=172445
X378 5 VIA1_C_CDNS_7194277470811 $T=214955 177475 0 0 $X=214035 $Y=177285
X379 5 VIA1_C_CDNS_7194277470811 $T=217155 59835 0 0 $X=216235 $Y=59645
X380 5 VIA1_C_CDNS_7194277470811 $T=217155 172635 0 0 $X=216235 $Y=172445
X381 5 VIA1_C_CDNS_7194277470811 $T=217155 177475 0 0 $X=216235 $Y=177285
X382 5 VIA1_C_CDNS_7194277470811 $T=221675 48755 0 0 $X=220755 $Y=48565
X383 7 VIA1_C_CDNS_7194277470811 $T=221675 54375 0 0 $X=220755 $Y=54185
X384 7 VIA1_C_CDNS_7194277470811 $T=221675 73175 0 0 $X=220755 $Y=72985
X385 7 VIA1_C_CDNS_7194277470811 $T=221675 91975 0 0 $X=220755 $Y=91785
X386 7 VIA1_C_CDNS_7194277470811 $T=221675 110775 0 0 $X=220755 $Y=110585
X387 7 VIA1_C_CDNS_7194277470811 $T=221675 129575 0 0 $X=220755 $Y=129385
X388 7 VIA1_C_CDNS_7194277470811 $T=221675 148375 0 0 $X=220755 $Y=148185
X389 5 VIA1_C_CDNS_7194277470811 $T=221675 172635 0 0 $X=220755 $Y=172445
X390 5 VIA1_C_CDNS_7194277470811 $T=226195 59835 0 0 $X=225275 $Y=59645
X391 14 VIA1_C_CDNS_7194277470811 $T=226195 77075 0 0 $X=225275 $Y=76885
X392 14 VIA1_C_CDNS_7194277470811 $T=226195 95875 0 0 $X=225275 $Y=95685
X393 14 VIA1_C_CDNS_7194277470811 $T=226195 133475 0 0 $X=225275 $Y=133285
X394 14 VIA1_C_CDNS_7194277470811 $T=226195 152275 0 0 $X=225275 $Y=152085
X395 14 VIA1_C_CDNS_7194277470811 $T=226195 171075 0 0 $X=225275 $Y=170885
X396 5 VIA1_C_CDNS_7194277470811 $T=226195 177475 0 0 $X=225275 $Y=177285
X397 5 VIA1_C_CDNS_7194277470811 $T=228395 59835 0 0 $X=227475 $Y=59645
X398 5 VIA1_C_CDNS_7194277470811 $T=228395 177475 0 0 $X=227475 $Y=177285
X399 5 VIA1_C_CDNS_7194277470811 $T=228965 172635 0 0 $X=228045 $Y=172445
X400 5 VIA1_C_CDNS_7194277470811 $T=232915 48755 0 0 $X=231995 $Y=48565
X401 7 VIA1_C_CDNS_7194277470811 $T=232915 54375 0 0 $X=231995 $Y=54185
X402 7 VIA1_C_CDNS_7194277470811 $T=232915 73175 0 0 $X=231995 $Y=72985
X403 7 VIA1_C_CDNS_7194277470811 $T=232915 91975 0 0 $X=231995 $Y=91785
X404 7 VIA1_C_CDNS_7194277470811 $T=232915 110775 0 0 $X=231995 $Y=110585
X405 7 VIA1_C_CDNS_7194277470811 $T=232915 129575 0 0 $X=231995 $Y=129385
X406 7 VIA1_C_CDNS_7194277470811 $T=232915 148375 0 0 $X=231995 $Y=148185
X407 5 VIA1_C_CDNS_7194277470811 $T=232915 172635 0 0 $X=231995 $Y=172445
X408 5 VIA1_C_CDNS_7194277470811 $T=237435 59835 0 0 $X=236515 $Y=59645
X409 15 VIA1_C_CDNS_7194277470811 $T=237435 76295 0 0 $X=236515 $Y=76105
X410 15 VIA1_C_CDNS_7194277470811 $T=237435 95095 0 0 $X=236515 $Y=94905
X411 15 VIA1_C_CDNS_7194277470811 $T=237435 132695 0 0 $X=236515 $Y=132505
X412 15 VIA1_C_CDNS_7194277470811 $T=237435 151495 0 0 $X=236515 $Y=151305
X413 14 VIA1_C_CDNS_7194277470811 $T=237435 171075 0 0 $X=236515 $Y=170885
X414 5 VIA1_C_CDNS_7194277470811 $T=237435 177475 0 0 $X=236515 $Y=177285
X415 5 VIA1_C_CDNS_7194277470811 $T=239635 59835 0 0 $X=238715 $Y=59645
X416 5 VIA1_C_CDNS_7194277470811 $T=239635 177475 0 0 $X=238715 $Y=177285
X417 5 VIA1_C_CDNS_7194277470811 $T=240205 172635 0 0 $X=239285 $Y=172445
X418 5 VIA1_C_CDNS_7194277470811 $T=244155 48755 0 0 $X=243235 $Y=48565
X419 7 VIA1_C_CDNS_7194277470811 $T=244155 54375 0 0 $X=243235 $Y=54185
X420 7 VIA1_C_CDNS_7194277470811 $T=244155 73175 0 0 $X=243235 $Y=72985
X421 7 VIA1_C_CDNS_7194277470811 $T=244155 91975 0 0 $X=243235 $Y=91785
X422 7 VIA1_C_CDNS_7194277470811 $T=244155 110775 0 0 $X=243235 $Y=110585
X423 7 VIA1_C_CDNS_7194277470811 $T=244155 129575 0 0 $X=243235 $Y=129385
X424 7 VIA1_C_CDNS_7194277470811 $T=244155 148375 0 0 $X=243235 $Y=148185
X425 5 VIA1_C_CDNS_7194277470811 $T=244155 172635 0 0 $X=243235 $Y=172445
X426 5 VIA1_C_CDNS_7194277470811 $T=248675 59835 0 0 $X=247755 $Y=59645
X427 15 VIA1_C_CDNS_7194277470811 $T=248675 76295 0 0 $X=247755 $Y=76105
X428 16 VIA1_C_CDNS_7194277470811 $T=248675 94315 0 0 $X=247755 $Y=94125
X429 16 VIA1_C_CDNS_7194277470811 $T=248675 131915 0 0 $X=247755 $Y=131725
X430 16 VIA1_C_CDNS_7194277470811 $T=248675 150715 0 0 $X=247755 $Y=150525
X431 14 VIA1_C_CDNS_7194277470811 $T=248675 171075 0 0 $X=247755 $Y=170885
X432 5 VIA1_C_CDNS_7194277470811 $T=248675 177475 0 0 $X=247755 $Y=177285
X433 5 VIA1_C_CDNS_7194277470811 $T=250875 59835 0 0 $X=249955 $Y=59645
X434 5 VIA1_C_CDNS_7194277470811 $T=250875 177475 0 0 $X=249955 $Y=177285
X435 5 VIA1_C_CDNS_7194277470811 $T=251445 172635 0 0 $X=250525 $Y=172445
X436 5 VIA1_C_CDNS_7194277470811 $T=255395 48755 0 0 $X=254475 $Y=48565
X437 7 VIA1_C_CDNS_7194277470811 $T=255395 54375 0 0 $X=254475 $Y=54185
X438 7 VIA1_C_CDNS_7194277470811 $T=255395 73175 0 0 $X=254475 $Y=72985
X439 7 VIA1_C_CDNS_7194277470811 $T=255395 91975 0 0 $X=254475 $Y=91785
X440 7 VIA1_C_CDNS_7194277470811 $T=255395 110775 0 0 $X=254475 $Y=110585
X441 7 VIA1_C_CDNS_7194277470811 $T=255395 129575 0 0 $X=254475 $Y=129385
X442 7 VIA1_C_CDNS_7194277470811 $T=255395 148375 0 0 $X=254475 $Y=148185
X443 5 VIA1_C_CDNS_7194277470811 $T=255395 172635 0 0 $X=254475 $Y=172445
X444 5 VIA1_C_CDNS_7194277470811 $T=259915 59835 0 0 $X=258995 $Y=59645
X445 15 VIA1_C_CDNS_7194277470811 $T=259915 76295 0 0 $X=258995 $Y=76105
X446 18 VIA1_C_CDNS_7194277470811 $T=259915 96655 0 0 $X=258995 $Y=96465
X447 18 VIA1_C_CDNS_7194277470811 $T=259915 134255 0 0 $X=258995 $Y=134065
X448 18 VIA1_C_CDNS_7194277470811 $T=259915 153055 0 0 $X=258995 $Y=152865
X449 14 VIA1_C_CDNS_7194277470811 $T=259915 171075 0 0 $X=258995 $Y=170885
X450 5 VIA1_C_CDNS_7194277470811 $T=259915 177475 0 0 $X=258995 $Y=177285
X451 5 VIA1_C_CDNS_7194277470811 $T=262115 59835 0 0 $X=261195 $Y=59645
X452 5 VIA1_C_CDNS_7194277470811 $T=262115 177475 0 0 $X=261195 $Y=177285
X453 5 VIA1_C_CDNS_7194277470811 $T=262685 172635 0 0 $X=261765 $Y=172445
X454 5 VIA1_C_CDNS_7194277470811 $T=266635 48755 0 0 $X=265715 $Y=48565
X455 7 VIA1_C_CDNS_7194277470811 $T=266635 54375 0 0 $X=265715 $Y=54185
X456 7 VIA1_C_CDNS_7194277470811 $T=266635 73175 0 0 $X=265715 $Y=72985
X457 7 VIA1_C_CDNS_7194277470811 $T=266635 91975 0 0 $X=265715 $Y=91785
X458 7 VIA1_C_CDNS_7194277470811 $T=266635 110775 0 0 $X=265715 $Y=110585
X459 7 VIA1_C_CDNS_7194277470811 $T=266635 129575 0 0 $X=265715 $Y=129385
X460 7 VIA1_C_CDNS_7194277470811 $T=266635 148375 0 0 $X=265715 $Y=148185
X461 5 VIA1_C_CDNS_7194277470811 $T=266635 172635 0 0 $X=265715 $Y=172445
X462 5 VIA1_C_CDNS_7194277470811 $T=271155 59835 0 0 $X=270235 $Y=59645
X463 15 VIA1_C_CDNS_7194277470811 $T=271155 76295 0 0 $X=270235 $Y=76105
X464 20 VIA1_C_CDNS_7194277470811 $T=271155 93535 0 0 $X=270235 $Y=93345
X465 17 VIA1_C_CDNS_7194277470811 $T=271155 130355 0 0 $X=270235 $Y=130165
X466 20 VIA1_C_CDNS_7194277470811 $T=271155 149935 0 0 $X=270235 $Y=149745
X467 14 VIA1_C_CDNS_7194277470811 $T=271155 171075 0 0 $X=270235 $Y=170885
X468 5 VIA1_C_CDNS_7194277470811 $T=271155 177475 0 0 $X=270235 $Y=177285
X469 5 VIA1_C_CDNS_7194277470811 $T=273355 59835 0 0 $X=272435 $Y=59645
X470 5 VIA1_C_CDNS_7194277470811 $T=273355 177475 0 0 $X=272435 $Y=177285
X471 5 VIA1_C_CDNS_7194277470811 $T=273925 172635 0 0 $X=273005 $Y=172445
X472 5 VIA1_C_CDNS_7194277470811 $T=277875 48755 0 0 $X=276955 $Y=48565
X473 7 VIA1_C_CDNS_7194277470811 $T=277875 54375 0 0 $X=276955 $Y=54185
X474 7 VIA1_C_CDNS_7194277470811 $T=277875 73175 0 0 $X=276955 $Y=72985
X475 7 VIA1_C_CDNS_7194277470811 $T=277875 91975 0 0 $X=276955 $Y=91785
X476 7 VIA1_C_CDNS_7194277470811 $T=277875 110775 0 0 $X=276955 $Y=110585
X477 7 VIA1_C_CDNS_7194277470811 $T=277875 129575 0 0 $X=276955 $Y=129385
X478 7 VIA1_C_CDNS_7194277470811 $T=277875 148375 0 0 $X=276955 $Y=148185
X479 5 VIA1_C_CDNS_7194277470811 $T=277875 172635 0 0 $X=276955 $Y=172445
X480 5 VIA1_C_CDNS_7194277470811 $T=282395 59835 0 0 $X=281475 $Y=59645
X481 18 VIA1_C_CDNS_7194277470811 $T=282395 77855 0 0 $X=281475 $Y=77665
X482 20 VIA1_C_CDNS_7194277470811 $T=282395 93535 0 0 $X=281475 $Y=93345
X483 18 VIA1_C_CDNS_7194277470811 $T=282395 134255 0 0 $X=281475 $Y=134065
X484 20 VIA1_C_CDNS_7194277470811 $T=282395 149935 0 0 $X=281475 $Y=149745
X485 15 VIA1_C_CDNS_7194277470811 $T=282395 170295 0 0 $X=281475 $Y=170105
X486 5 VIA1_C_CDNS_7194277470811 $T=282395 177475 0 0 $X=281475 $Y=177285
X487 5 VIA1_C_CDNS_7194277470811 $T=284595 59835 0 0 $X=283675 $Y=59645
X488 5 VIA1_C_CDNS_7194277470811 $T=284595 177475 0 0 $X=283675 $Y=177285
X489 5 VIA1_C_CDNS_7194277470811 $T=285165 172635 0 0 $X=284245 $Y=172445
X490 5 VIA1_C_CDNS_7194277470811 $T=289115 48755 0 0 $X=288195 $Y=48565
X491 7 VIA1_C_CDNS_7194277470811 $T=289115 54375 0 0 $X=288195 $Y=54185
X492 7 VIA1_C_CDNS_7194277470811 $T=289115 73175 0 0 $X=288195 $Y=72985
X493 7 VIA1_C_CDNS_7194277470811 $T=289115 91975 0 0 $X=288195 $Y=91785
X494 7 VIA1_C_CDNS_7194277470811 $T=289115 110775 0 0 $X=288195 $Y=110585
X495 7 VIA1_C_CDNS_7194277470811 $T=289115 129575 0 0 $X=288195 $Y=129385
X496 7 VIA1_C_CDNS_7194277470811 $T=289115 148375 0 0 $X=288195 $Y=148185
X497 5 VIA1_C_CDNS_7194277470811 $T=289115 172635 0 0 $X=288195 $Y=172445
X498 5 VIA1_C_CDNS_7194277470811 $T=293635 59835 0 0 $X=292715 $Y=59645
X499 14 VIA1_C_CDNS_7194277470811 $T=293635 77075 0 0 $X=292715 $Y=76885
X500 18 VIA1_C_CDNS_7194277470811 $T=293635 96655 0 0 $X=292715 $Y=96465
X501 16 VIA1_C_CDNS_7194277470811 $T=293635 131915 0 0 $X=292715 $Y=131725
X502 18 VIA1_C_CDNS_7194277470811 $T=293635 153055 0 0 $X=292715 $Y=152865
X503 15 VIA1_C_CDNS_7194277470811 $T=293635 170295 0 0 $X=292715 $Y=170105
X504 5 VIA1_C_CDNS_7194277470811 $T=293635 177475 0 0 $X=292715 $Y=177285
X505 5 VIA1_C_CDNS_7194277470811 $T=295835 59835 0 0 $X=294915 $Y=59645
X506 5 VIA1_C_CDNS_7194277470811 $T=295835 177475 0 0 $X=294915 $Y=177285
X507 5 VIA1_C_CDNS_7194277470811 $T=296405 172635 0 0 $X=295485 $Y=172445
X508 5 VIA1_C_CDNS_7194277470811 $T=300355 48755 0 0 $X=299435 $Y=48565
X509 7 VIA1_C_CDNS_7194277470811 $T=300355 54375 0 0 $X=299435 $Y=54185
X510 7 VIA1_C_CDNS_7194277470811 $T=300355 73175 0 0 $X=299435 $Y=72985
X511 7 VIA1_C_CDNS_7194277470811 $T=300355 91975 0 0 $X=299435 $Y=91785
X512 7 VIA1_C_CDNS_7194277470811 $T=300355 110775 0 0 $X=299435 $Y=110585
X513 7 VIA1_C_CDNS_7194277470811 $T=300355 129575 0 0 $X=299435 $Y=129385
X514 7 VIA1_C_CDNS_7194277470811 $T=300355 148375 0 0 $X=299435 $Y=148185
X515 5 VIA1_C_CDNS_7194277470811 $T=300355 172635 0 0 $X=299435 $Y=172445
X516 5 VIA1_C_CDNS_7194277470811 $T=304875 59835 0 0 $X=303955 $Y=59645
X517 14 VIA1_C_CDNS_7194277470811 $T=304875 77075 0 0 $X=303955 $Y=76885
X518 16 VIA1_C_CDNS_7194277470811 $T=304875 94315 0 0 $X=303955 $Y=94125
X519 15 VIA1_C_CDNS_7194277470811 $T=304875 132695 0 0 $X=303955 $Y=132505
X520 16 VIA1_C_CDNS_7194277470811 $T=304875 150715 0 0 $X=303955 $Y=150525
X521 15 VIA1_C_CDNS_7194277470811 $T=304875 170295 0 0 $X=303955 $Y=170105
X522 5 VIA1_C_CDNS_7194277470811 $T=304875 177475 0 0 $X=303955 $Y=177285
X523 5 VIA1_C_CDNS_7194277470811 $T=307075 59835 0 0 $X=306155 $Y=59645
X524 5 VIA1_C_CDNS_7194277470811 $T=307075 177475 0 0 $X=306155 $Y=177285
X525 5 VIA1_C_CDNS_7194277470811 $T=307645 172635 0 0 $X=306725 $Y=172445
X526 5 VIA1_C_CDNS_7194277470811 $T=311595 48755 0 0 $X=310675 $Y=48565
X527 5 VIA1_C_CDNS_7194277470811 $T=311595 59835 0 0 $X=310675 $Y=59645
X528 7 VIA1_C_CDNS_7194277470811 $T=311595 73175 0 0 $X=310675 $Y=72985
X529 7 VIA1_C_CDNS_7194277470811 $T=311595 91975 0 0 $X=310675 $Y=91785
X530 7 VIA1_C_CDNS_7194277470811 $T=311595 110775 0 0 $X=310675 $Y=110585
X531 7 VIA1_C_CDNS_7194277470811 $T=311595 129575 0 0 $X=310675 $Y=129385
X532 7 VIA1_C_CDNS_7194277470811 $T=311595 148375 0 0 $X=310675 $Y=148185
X533 5 VIA1_C_CDNS_7194277470811 $T=311595 172635 0 0 $X=310675 $Y=172445
X534 5 VIA1_C_CDNS_7194277470811 $T=316115 59835 0 0 $X=315195 $Y=59645
X535 5 VIA1_C_CDNS_7194277470811 $T=316115 78635 0 0 $X=315195 $Y=78445
X536 15 VIA1_C_CDNS_7194277470811 $T=316115 95095 0 0 $X=315195 $Y=94905
X537 15 VIA1_C_CDNS_7194277470811 $T=316115 132695 0 0 $X=315195 $Y=132505
X538 15 VIA1_C_CDNS_7194277470811 $T=316115 151495 0 0 $X=315195 $Y=151305
X539 18 VIA1_C_CDNS_7194277470811 $T=316115 171855 0 0 $X=315195 $Y=171665
X540 5 VIA1_C_CDNS_7194277470811 $T=316115 177475 0 0 $X=315195 $Y=177285
X541 5 VIA1_C_CDNS_7194277470811 $T=318315 59835 0 0 $X=317395 $Y=59645
X542 5 VIA1_C_CDNS_7194277470811 $T=318315 177475 0 0 $X=317395 $Y=177285
X543 5 VIA1_C_CDNS_7194277470811 $T=318885 172635 0 0 $X=317965 $Y=172445
X544 5 VIA1_C_CDNS_7194277470811 $T=322835 48755 0 0 $X=321915 $Y=48565
X545 5 VIA1_C_CDNS_7194277470811 $T=322835 59835 0 0 $X=321915 $Y=59645
X546 7 VIA1_C_CDNS_7194277470811 $T=322835 73175 0 0 $X=321915 $Y=72985
X547 7 VIA1_C_CDNS_7194277470811 $T=322835 91975 0 0 $X=321915 $Y=91785
X548 7 VIA1_C_CDNS_7194277470811 $T=322835 110775 0 0 $X=321915 $Y=110585
X549 7 VIA1_C_CDNS_7194277470811 $T=322835 129575 0 0 $X=321915 $Y=129385
X550 7 VIA1_C_CDNS_7194277470811 $T=322835 148375 0 0 $X=321915 $Y=148185
X551 5 VIA1_C_CDNS_7194277470811 $T=322835 172635 0 0 $X=321915 $Y=172445
X552 5 VIA1_C_CDNS_7194277470811 $T=327355 59835 0 0 $X=326435 $Y=59645
X553 5 VIA1_C_CDNS_7194277470811 $T=327355 78635 0 0 $X=326435 $Y=78445
X554 14 VIA1_C_CDNS_7194277470811 $T=327355 95875 0 0 $X=326435 $Y=95685
X555 14 VIA1_C_CDNS_7194277470811 $T=327355 133475 0 0 $X=326435 $Y=133285
X556 14 VIA1_C_CDNS_7194277470811 $T=327355 152275 0 0 $X=326435 $Y=152085
X557 14 VIA1_C_CDNS_7194277470811 $T=327355 171075 0 0 $X=326435 $Y=170885
X558 5 VIA1_C_CDNS_7194277470811 $T=327355 177475 0 0 $X=326435 $Y=177285
X559 5 VIA1_C_CDNS_7194277470811 $T=329555 59835 0 0 $X=328635 $Y=59645
X560 5 VIA1_C_CDNS_7194277470811 $T=329555 177475 0 0 $X=328635 $Y=177285
X561 5 VIA1_C_CDNS_7194277470811 $T=330125 172635 0 0 $X=329205 $Y=172445
X562 5 VIA1_C_CDNS_7194277470811 $T=334075 48755 0 0 $X=333155 $Y=48565
X563 5 VIA1_C_CDNS_7194277470811 $T=334075 59835 0 0 $X=333155 $Y=59645
X564 7 VIA1_C_CDNS_7194277470811 $T=334075 73175 0 0 $X=333155 $Y=72985
X565 7 VIA1_C_CDNS_7194277470811 $T=334075 91975 0 0 $X=333155 $Y=91785
X566 7 VIA1_C_CDNS_7194277470811 $T=334075 110775 0 0 $X=333155 $Y=110585
X567 7 VIA1_C_CDNS_7194277470811 $T=334075 129575 0 0 $X=333155 $Y=129385
X568 7 VIA1_C_CDNS_7194277470811 $T=334075 148375 0 0 $X=333155 $Y=148185
X569 5 VIA1_C_CDNS_7194277470811 $T=334075 172635 0 0 $X=333155 $Y=172445
X570 5 VIA1_C_CDNS_7194277470811 $T=338595 59835 0 0 $X=337675 $Y=59645
X571 5 VIA1_C_CDNS_7194277470811 $T=338595 78635 0 0 $X=337675 $Y=78445
X572 14 VIA1_C_CDNS_7194277470811 $T=338595 95875 0 0 $X=337675 $Y=95685
X573 14 VIA1_C_CDNS_7194277470811 $T=338595 133475 0 0 $X=337675 $Y=133285
X574 14 VIA1_C_CDNS_7194277470811 $T=338595 152275 0 0 $X=337675 $Y=152085
X575 14 VIA1_C_CDNS_7194277470811 $T=338595 171075 0 0 $X=337675 $Y=170885
X576 5 VIA1_C_CDNS_7194277470811 $T=338595 177475 0 0 $X=337675 $Y=177285
X577 5 VIA1_C_CDNS_7194277470811 $T=340795 59835 0 0 $X=339875 $Y=59645
X578 5 VIA1_C_CDNS_7194277470811 $T=340795 177475 0 0 $X=339875 $Y=177285
X579 5 VIA1_C_CDNS_7194277470811 $T=341365 172635 0 0 $X=340445 $Y=172445
X580 5 VIA1_C_CDNS_7194277470811 $T=345315 48755 0 0 $X=344395 $Y=48565
X581 5 VIA1_C_CDNS_7194277470811 $T=345315 59835 0 0 $X=344395 $Y=59645
X582 7 VIA1_C_CDNS_7194277470811 $T=345315 73175 0 0 $X=344395 $Y=72985
X583 7 VIA1_C_CDNS_7194277470811 $T=345315 91975 0 0 $X=344395 $Y=91785
X584 7 VIA1_C_CDNS_7194277470811 $T=345315 110775 0 0 $X=344395 $Y=110585
X585 7 VIA1_C_CDNS_7194277470811 $T=345315 129575 0 0 $X=344395 $Y=129385
X586 7 VIA1_C_CDNS_7194277470811 $T=345315 148375 0 0 $X=344395 $Y=148185
X587 5 VIA1_C_CDNS_7194277470811 $T=345315 172635 0 0 $X=344395 $Y=172445
X588 5 VIA1_C_CDNS_7194277470811 $T=349835 59835 0 0 $X=348915 $Y=59645
X589 5 VIA1_C_CDNS_7194277470811 $T=349835 78635 0 0 $X=348915 $Y=78445
X590 14 VIA1_C_CDNS_7194277470811 $T=349835 95875 0 0 $X=348915 $Y=95685
X591 14 VIA1_C_CDNS_7194277470811 $T=349835 133475 0 0 $X=348915 $Y=133285
X592 14 VIA1_C_CDNS_7194277470811 $T=349835 152275 0 0 $X=348915 $Y=152085
X593 14 VIA1_C_CDNS_7194277470811 $T=349835 171075 0 0 $X=348915 $Y=170885
X594 5 VIA1_C_CDNS_7194277470811 $T=349835 177475 0 0 $X=348915 $Y=177285
X595 5 VIA1_C_CDNS_7194277470811 $T=352035 59835 0 0 $X=351115 $Y=59645
X596 5 VIA1_C_CDNS_7194277470811 $T=352035 177475 0 0 $X=351115 $Y=177285
X597 5 VIA1_C_CDNS_7194277470811 $T=352605 172635 0 0 $X=351685 $Y=172445
X598 5 VIA1_C_CDNS_7194277470811 $T=356555 48755 0 0 $X=355635 $Y=48565
X599 5 VIA1_C_CDNS_7194277470811 $T=356555 59835 0 0 $X=355635 $Y=59645
X600 7 VIA1_C_CDNS_7194277470811 $T=356555 73175 0 0 $X=355635 $Y=72985
X601 7 VIA1_C_CDNS_7194277470811 $T=356555 91975 0 0 $X=355635 $Y=91785
X602 7 VIA1_C_CDNS_7194277470811 $T=356555 110775 0 0 $X=355635 $Y=110585
X603 7 VIA1_C_CDNS_7194277470811 $T=356555 129575 0 0 $X=355635 $Y=129385
X604 7 VIA1_C_CDNS_7194277470811 $T=356555 148375 0 0 $X=355635 $Y=148185
X605 5 VIA1_C_CDNS_7194277470811 $T=356555 172635 0 0 $X=355635 $Y=172445
X606 5 VIA1_C_CDNS_7194277470811 $T=361075 59835 0 0 $X=360155 $Y=59645
X607 5 VIA1_C_CDNS_7194277470811 $T=361075 78635 0 0 $X=360155 $Y=78445
X608 14 VIA1_C_CDNS_7194277470811 $T=361075 95875 0 0 $X=360155 $Y=95685
X609 14 VIA1_C_CDNS_7194277470811 $T=361075 133475 0 0 $X=360155 $Y=133285
X610 14 VIA1_C_CDNS_7194277470811 $T=361075 152275 0 0 $X=360155 $Y=152085
X611 14 VIA1_C_CDNS_7194277470811 $T=361075 171075 0 0 $X=360155 $Y=170885
X612 5 VIA1_C_CDNS_7194277470811 $T=361075 177475 0 0 $X=360155 $Y=177285
X613 5 VIA1_C_CDNS_7194277470811 $T=363275 59835 0 0 $X=362355 $Y=59645
X614 5 VIA1_C_CDNS_7194277470811 $T=363275 177475 0 0 $X=362355 $Y=177285
X615 5 VIA1_C_CDNS_7194277470811 $T=363845 172635 0 0 $X=362925 $Y=172445
X616 5 VIA1_C_CDNS_7194277470811 $T=367795 48755 0 0 $X=366875 $Y=48565
X617 5 VIA1_C_CDNS_7194277470811 $T=367795 59835 0 0 $X=366875 $Y=59645
X618 5 VIA1_C_CDNS_7194277470811 $T=367795 78635 0 0 $X=366875 $Y=78445
X619 5 VIA1_C_CDNS_7194277470811 $T=367795 97435 0 0 $X=366875 $Y=97245
X620 5 VIA1_C_CDNS_7194277470811 $T=367795 116235 0 0 $X=366875 $Y=116045
X621 5 VIA1_C_CDNS_7194277470811 $T=367795 135035 0 0 $X=366875 $Y=134845
X622 5 VIA1_C_CDNS_7194277470811 $T=367795 153835 0 0 $X=366875 $Y=153645
X623 5 VIA1_C_CDNS_7194277470811 $T=367795 172635 0 0 $X=366875 $Y=172445
X624 5 VIA1_C_CDNS_7194277470811 $T=373065 59835 0 0 $X=372145 $Y=59645
X625 5 VIA1_C_CDNS_7194277470811 $T=373065 78635 0 0 $X=372145 $Y=78445
X626 5 VIA1_C_CDNS_7194277470811 $T=373065 97435 0 0 $X=372145 $Y=97245
X627 5 VIA1_C_CDNS_7194277470811 $T=373065 116235 0 0 $X=372145 $Y=116045
X628 5 VIA1_C_CDNS_7194277470811 $T=373065 135035 0 0 $X=372145 $Y=134845
X629 5 VIA1_C_CDNS_7194277470811 $T=373065 153835 0 0 $X=372145 $Y=153645
X630 5 VIA1_C_CDNS_7194277470811 $T=373065 172635 0 0 $X=372145 $Y=172445
X631 5 VIA1_C_CDNS_7194277470811 $T=373065 177475 0 0 $X=372145 $Y=177285
X632 19 VIA2_C_CDNS_7194277470812 $T=184405 53595 0 0 $X=183485 $Y=53405
X633 19 VIA2_C_CDNS_7194277470812 $T=184405 72395 0 0 $X=183485 $Y=72205
X634 19 VIA2_C_CDNS_7194277470812 $T=184405 91195 0 0 $X=183485 $Y=91005
X635 19 VIA2_C_CDNS_7194277470812 $T=184405 109995 0 0 $X=183485 $Y=109805
X636 19 VIA2_C_CDNS_7194277470812 $T=184405 128795 0 0 $X=183485 $Y=128605
X637 19 VIA2_C_CDNS_7194277470812 $T=184405 147595 0 0 $X=183485 $Y=147405
X638 19 VIA2_C_CDNS_7194277470812 $T=184405 166395 0 0 $X=183485 $Y=166205
X639 7 VIA2_C_CDNS_7194277470812 $T=186685 54375 0 0 $X=185765 $Y=54185
X640 7 VIA2_C_CDNS_7194277470812 $T=186685 73175 0 0 $X=185765 $Y=72985
X641 7 VIA2_C_CDNS_7194277470812 $T=186685 91975 0 0 $X=185765 $Y=91785
X642 7 VIA2_C_CDNS_7194277470812 $T=186685 110775 0 0 $X=185765 $Y=110585
X643 7 VIA2_C_CDNS_7194277470812 $T=186685 129575 0 0 $X=185765 $Y=129385
X644 7 VIA2_C_CDNS_7194277470812 $T=186685 148375 0 0 $X=185765 $Y=148185
X645 7 VIA2_C_CDNS_7194277470812 $T=186685 167175 0 0 $X=185765 $Y=166985
X646 17 VIA2_C_CDNS_7194277470812 $T=188965 55155 0 0 $X=188045 $Y=54965
X647 17 VIA2_C_CDNS_7194277470812 $T=188965 73955 0 0 $X=188045 $Y=73765
X648 17 VIA2_C_CDNS_7194277470812 $T=188965 92755 0 0 $X=188045 $Y=92565
X649 17 VIA2_C_CDNS_7194277470812 $T=188965 111555 0 0 $X=188045 $Y=111365
X650 17 VIA2_C_CDNS_7194277470812 $T=188965 130355 0 0 $X=188045 $Y=130165
X651 17 VIA2_C_CDNS_7194277470812 $T=188965 149155 0 0 $X=188045 $Y=148965
X652 17 VIA2_C_CDNS_7194277470812 $T=188965 167955 0 0 $X=188045 $Y=167765
X653 20 VIA2_C_CDNS_7194277470812 $T=191245 55935 0 0 $X=190325 $Y=55745
X654 20 VIA2_C_CDNS_7194277470812 $T=191245 74735 0 0 $X=190325 $Y=74545
X655 20 VIA2_C_CDNS_7194277470812 $T=191245 93535 0 0 $X=190325 $Y=93345
X656 20 VIA2_C_CDNS_7194277470812 $T=191245 112335 0 0 $X=190325 $Y=112145
X657 20 VIA2_C_CDNS_7194277470812 $T=191245 131135 0 0 $X=190325 $Y=130945
X658 20 VIA2_C_CDNS_7194277470812 $T=191245 149935 0 0 $X=190325 $Y=149745
X659 20 VIA2_C_CDNS_7194277470812 $T=191245 168735 0 0 $X=190325 $Y=168545
X660 16 VIA2_C_CDNS_7194277470812 $T=193525 56715 0 0 $X=192605 $Y=56525
X661 16 VIA2_C_CDNS_7194277470812 $T=193525 75515 0 0 $X=192605 $Y=75325
X662 16 VIA2_C_CDNS_7194277470812 $T=193525 94315 0 0 $X=192605 $Y=94125
X663 16 VIA2_C_CDNS_7194277470812 $T=193525 113115 0 0 $X=192605 $Y=112925
X664 16 VIA2_C_CDNS_7194277470812 $T=193525 131915 0 0 $X=192605 $Y=131725
X665 16 VIA2_C_CDNS_7194277470812 $T=193525 150715 0 0 $X=192605 $Y=150525
X666 16 VIA2_C_CDNS_7194277470812 $T=193525 169515 0 0 $X=192605 $Y=169325
X667 15 VIA2_C_CDNS_7194277470812 $T=195805 57495 0 0 $X=194885 $Y=57305
X668 15 VIA2_C_CDNS_7194277470812 $T=195805 76295 0 0 $X=194885 $Y=76105
X669 15 VIA2_C_CDNS_7194277470812 $T=195805 95095 0 0 $X=194885 $Y=94905
X670 15 VIA2_C_CDNS_7194277470812 $T=195805 113895 0 0 $X=194885 $Y=113705
X671 15 VIA2_C_CDNS_7194277470812 $T=195805 132695 0 0 $X=194885 $Y=132505
X672 15 VIA2_C_CDNS_7194277470812 $T=195805 151495 0 0 $X=194885 $Y=151305
X673 15 VIA2_C_CDNS_7194277470812 $T=195805 170295 0 0 $X=194885 $Y=170105
X674 14 VIA2_C_CDNS_7194277470812 $T=198085 58275 0 0 $X=197165 $Y=58085
X675 14 VIA2_C_CDNS_7194277470812 $T=198085 77075 0 0 $X=197165 $Y=76885
X676 14 VIA2_C_CDNS_7194277470812 $T=198085 95875 0 0 $X=197165 $Y=95685
X677 14 VIA2_C_CDNS_7194277470812 $T=198085 114675 0 0 $X=197165 $Y=114485
X678 14 VIA2_C_CDNS_7194277470812 $T=198085 133475 0 0 $X=197165 $Y=133285
X679 14 VIA2_C_CDNS_7194277470812 $T=198085 152275 0 0 $X=197165 $Y=152085
X680 14 VIA2_C_CDNS_7194277470812 $T=198085 171075 0 0 $X=197165 $Y=170885
X681 18 VIA2_C_CDNS_7194277470812 $T=200365 59055 0 0 $X=199445 $Y=58865
X682 18 VIA2_C_CDNS_7194277470812 $T=200365 77855 0 0 $X=199445 $Y=77665
X683 18 VIA2_C_CDNS_7194277470812 $T=200365 96655 0 0 $X=199445 $Y=96465
X684 18 VIA2_C_CDNS_7194277470812 $T=200365 115455 0 0 $X=199445 $Y=115265
X685 18 VIA2_C_CDNS_7194277470812 $T=200365 134255 0 0 $X=199445 $Y=134065
X686 18 VIA2_C_CDNS_7194277470812 $T=200365 153055 0 0 $X=199445 $Y=152865
X687 18 VIA2_C_CDNS_7194277470812 $T=200365 171855 0 0 $X=199445 $Y=171665
X688 5 VIA2_C_CDNS_7194277470812 $T=202645 48755 0 0 $X=201725 $Y=48565
X689 5 VIA2_C_CDNS_7194277470812 $T=202645 59835 0 0 $X=201725 $Y=59645
X690 5 VIA2_C_CDNS_7194277470812 $T=202645 78635 0 0 $X=201725 $Y=78445
X691 5 VIA2_C_CDNS_7194277470812 $T=202645 97435 0 0 $X=201725 $Y=97245
X692 5 VIA2_C_CDNS_7194277470812 $T=202645 116235 0 0 $X=201725 $Y=116045
X693 5 VIA2_C_CDNS_7194277470812 $T=202645 135035 0 0 $X=201725 $Y=134845
X694 5 VIA2_C_CDNS_7194277470812 $T=202645 153835 0 0 $X=201725 $Y=153645
X695 5 VIA2_C_CDNS_7194277470812 $T=202645 172635 0 0 $X=201725 $Y=172445
X696 5 VIA2_C_CDNS_7194277470812 $T=202645 177475 0 0 $X=201725 $Y=177285
X697 5 VIA2_C_CDNS_7194277470812 $T=375585 48755 0 0 $X=374665 $Y=48565
X698 5 VIA2_C_CDNS_7194277470812 $T=375585 59835 0 0 $X=374665 $Y=59645
X699 5 VIA2_C_CDNS_7194277470812 $T=375585 78635 0 0 $X=374665 $Y=78445
X700 5 VIA2_C_CDNS_7194277470812 $T=375585 97435 0 0 $X=374665 $Y=97245
X701 5 VIA2_C_CDNS_7194277470812 $T=375585 116235 0 0 $X=374665 $Y=116045
X702 5 VIA2_C_CDNS_7194277470812 $T=375585 135035 0 0 $X=374665 $Y=134845
X703 5 VIA2_C_CDNS_7194277470812 $T=375585 153835 0 0 $X=374665 $Y=153645
X704 5 VIA2_C_CDNS_7194277470812 $T=375585 172635 0 0 $X=374665 $Y=172445
X705 5 VIA2_C_CDNS_7194277470812 $T=375585 177475 0 0 $X=374665 $Y=177285
X706 19 VIA2_C_CDNS_7194277470812 $T=377865 53595 0 0 $X=376945 $Y=53405
X707 19 VIA2_C_CDNS_7194277470812 $T=377865 72395 0 0 $X=376945 $Y=72205
X708 19 VIA2_C_CDNS_7194277470812 $T=377865 91195 0 0 $X=376945 $Y=91005
X709 19 VIA2_C_CDNS_7194277470812 $T=377865 109995 0 0 $X=376945 $Y=109805
X710 19 VIA2_C_CDNS_7194277470812 $T=377865 128795 0 0 $X=376945 $Y=128605
X711 19 VIA2_C_CDNS_7194277470812 $T=377865 147595 0 0 $X=376945 $Y=147405
X712 19 VIA2_C_CDNS_7194277470812 $T=377865 166395 0 0 $X=376945 $Y=166205
X713 7 VIA2_C_CDNS_7194277470812 $T=380145 54375 0 0 $X=379225 $Y=54185
X714 7 VIA2_C_CDNS_7194277470812 $T=380145 73175 0 0 $X=379225 $Y=72985
X715 7 VIA2_C_CDNS_7194277470812 $T=380145 91975 0 0 $X=379225 $Y=91785
X716 7 VIA2_C_CDNS_7194277470812 $T=380145 110775 0 0 $X=379225 $Y=110585
X717 7 VIA2_C_CDNS_7194277470812 $T=380145 129575 0 0 $X=379225 $Y=129385
X718 7 VIA2_C_CDNS_7194277470812 $T=380145 148375 0 0 $X=379225 $Y=148185
X719 7 VIA2_C_CDNS_7194277470812 $T=380145 167175 0 0 $X=379225 $Y=166985
X720 17 VIA2_C_CDNS_7194277470812 $T=382425 55155 0 0 $X=381505 $Y=54965
X721 17 VIA2_C_CDNS_7194277470812 $T=382425 73955 0 0 $X=381505 $Y=73765
X722 17 VIA2_C_CDNS_7194277470812 $T=382425 92755 0 0 $X=381505 $Y=92565
X723 17 VIA2_C_CDNS_7194277470812 $T=382425 111555 0 0 $X=381505 $Y=111365
X724 17 VIA2_C_CDNS_7194277470812 $T=382425 130355 0 0 $X=381505 $Y=130165
X725 17 VIA2_C_CDNS_7194277470812 $T=382425 149155 0 0 $X=381505 $Y=148965
X726 17 VIA2_C_CDNS_7194277470812 $T=382425 167955 0 0 $X=381505 $Y=167765
X727 20 VIA2_C_CDNS_7194277470812 $T=384705 55935 0 0 $X=383785 $Y=55745
X728 20 VIA2_C_CDNS_7194277470812 $T=384705 74735 0 0 $X=383785 $Y=74545
X729 20 VIA2_C_CDNS_7194277470812 $T=384705 93535 0 0 $X=383785 $Y=93345
X730 20 VIA2_C_CDNS_7194277470812 $T=384705 112335 0 0 $X=383785 $Y=112145
X731 20 VIA2_C_CDNS_7194277470812 $T=384705 131135 0 0 $X=383785 $Y=130945
X732 20 VIA2_C_CDNS_7194277470812 $T=384705 149935 0 0 $X=383785 $Y=149745
X733 20 VIA2_C_CDNS_7194277470812 $T=384705 168735 0 0 $X=383785 $Y=168545
X734 16 VIA2_C_CDNS_7194277470812 $T=386985 56715 0 0 $X=386065 $Y=56525
X735 16 VIA2_C_CDNS_7194277470812 $T=386985 75515 0 0 $X=386065 $Y=75325
X736 16 VIA2_C_CDNS_7194277470812 $T=386985 94315 0 0 $X=386065 $Y=94125
X737 16 VIA2_C_CDNS_7194277470812 $T=386985 113115 0 0 $X=386065 $Y=112925
X738 16 VIA2_C_CDNS_7194277470812 $T=386985 131915 0 0 $X=386065 $Y=131725
X739 16 VIA2_C_CDNS_7194277470812 $T=386985 150715 0 0 $X=386065 $Y=150525
X740 16 VIA2_C_CDNS_7194277470812 $T=386985 169515 0 0 $X=386065 $Y=169325
X741 15 VIA2_C_CDNS_7194277470812 $T=389265 57495 0 0 $X=388345 $Y=57305
X742 15 VIA2_C_CDNS_7194277470812 $T=389265 76295 0 0 $X=388345 $Y=76105
X743 15 VIA2_C_CDNS_7194277470812 $T=389265 95095 0 0 $X=388345 $Y=94905
X744 15 VIA2_C_CDNS_7194277470812 $T=389265 113895 0 0 $X=388345 $Y=113705
X745 15 VIA2_C_CDNS_7194277470812 $T=389265 132695 0 0 $X=388345 $Y=132505
X746 15 VIA2_C_CDNS_7194277470812 $T=389265 151495 0 0 $X=388345 $Y=151305
X747 15 VIA2_C_CDNS_7194277470812 $T=389265 170295 0 0 $X=388345 $Y=170105
X748 14 VIA2_C_CDNS_7194277470812 $T=391545 58275 0 0 $X=390625 $Y=58085
X749 14 VIA2_C_CDNS_7194277470812 $T=391545 77075 0 0 $X=390625 $Y=76885
X750 14 VIA2_C_CDNS_7194277470812 $T=391545 95875 0 0 $X=390625 $Y=95685
X751 14 VIA2_C_CDNS_7194277470812 $T=391545 114675 0 0 $X=390625 $Y=114485
X752 14 VIA2_C_CDNS_7194277470812 $T=391545 133475 0 0 $X=390625 $Y=133285
X753 14 VIA2_C_CDNS_7194277470812 $T=391545 152275 0 0 $X=390625 $Y=152085
X754 14 VIA2_C_CDNS_7194277470812 $T=391545 171075 0 0 $X=390625 $Y=170885
X755 18 VIA2_C_CDNS_7194277470812 $T=393825 59055 0 0 $X=392905 $Y=58865
X756 18 VIA2_C_CDNS_7194277470812 $T=393825 77855 0 0 $X=392905 $Y=77665
X757 18 VIA2_C_CDNS_7194277470812 $T=393825 96655 0 0 $X=392905 $Y=96465
X758 18 VIA2_C_CDNS_7194277470812 $T=393825 115455 0 0 $X=392905 $Y=115265
X759 18 VIA2_C_CDNS_7194277470812 $T=393825 134255 0 0 $X=392905 $Y=134065
X760 18 VIA2_C_CDNS_7194277470812 $T=393825 153055 0 0 $X=392905 $Y=152865
X761 18 VIA2_C_CDNS_7194277470812 $T=393825 171855 0 0 $X=392905 $Y=171665
X762 18 VIA1_C_CDNS_7194277470813 $T=223665 38490 1 0 $X=223265 $Y=37520
X763 21 VIA1_C_CDNS_7194277470813 $T=225205 40770 1 0 $X=224805 $Y=39800
X764 18 VIA1_C_CDNS_7194277470813 $T=226745 38490 1 0 $X=226345 $Y=37520
X765 21 VIA1_C_CDNS_7194277470813 $T=228285 40770 1 0 $X=227885 $Y=39800
X766 18 VIA1_C_CDNS_7194277470813 $T=229825 38490 1 0 $X=229425 $Y=37520
X767 21 VIA1_C_CDNS_7194277470813 $T=231365 40770 1 0 $X=230965 $Y=39800
X768 18 VIA1_C_CDNS_7194277470813 $T=232905 38490 1 0 $X=232505 $Y=37520
X769 21 VIA1_C_CDNS_7194277470813 $T=234445 40770 1 0 $X=234045 $Y=39800
X770 18 VIA1_C_CDNS_7194277470813 $T=235985 38490 1 0 $X=235585 $Y=37520
X771 21 VIA1_C_CDNS_7194277470813 $T=237525 40770 1 0 $X=237125 $Y=39800
X772 18 VIA1_C_CDNS_7194277470813 $T=239065 38490 1 0 $X=238665 $Y=37520
X773 14 VIA1_C_CDNS_7194277470813 $T=246485 40770 1 0 $X=246085 $Y=39800
X774 22 VIA1_C_CDNS_7194277470813 $T=248025 38490 1 0 $X=247625 $Y=37520
X775 14 VIA1_C_CDNS_7194277470813 $T=249565 40770 1 0 $X=249165 $Y=39800
X776 22 VIA1_C_CDNS_7194277470813 $T=251105 38490 1 0 $X=250705 $Y=37520
X777 14 VIA1_C_CDNS_7194277470813 $T=252645 40770 1 0 $X=252245 $Y=39800
X778 22 VIA1_C_CDNS_7194277470813 $T=254185 38490 1 0 $X=253785 $Y=37520
X779 14 VIA1_C_CDNS_7194277470813 $T=255725 40770 1 0 $X=255325 $Y=39800
X780 22 VIA1_C_CDNS_7194277470813 $T=257265 38490 1 0 $X=256865 $Y=37520
X781 14 VIA1_C_CDNS_7194277470813 $T=258805 40770 1 0 $X=258405 $Y=39800
X782 22 VIA1_C_CDNS_7194277470813 $T=260345 38490 1 0 $X=259945 $Y=37520
X783 14 VIA1_C_CDNS_7194277470813 $T=261885 40770 1 0 $X=261485 $Y=39800
X784 22 VIA1_C_CDNS_7194277470813 $T=263425 38490 1 0 $X=263025 $Y=37520
X785 14 VIA1_C_CDNS_7194277470813 $T=264965 40770 1 0 $X=264565 $Y=39800
X786 22 VIA1_C_CDNS_7194277470813 $T=266505 38490 1 0 $X=266105 $Y=37520
X787 14 VIA1_C_CDNS_7194277470813 $T=268045 40770 1 0 $X=267645 $Y=39800
X788 22 VIA1_C_CDNS_7194277470813 $T=269585 38490 1 0 $X=269185 $Y=37520
X789 14 VIA1_C_CDNS_7194277470813 $T=271125 40770 1 0 $X=270725 $Y=39800
X790 22 VIA1_C_CDNS_7194277470813 $T=272665 38490 1 0 $X=272265 $Y=37520
X791 14 VIA1_C_CDNS_7194277470813 $T=274205 40770 1 0 $X=273805 $Y=39800
X792 22 VIA1_C_CDNS_7194277470813 $T=275745 38490 1 0 $X=275345 $Y=37520
X793 14 VIA1_C_CDNS_7194277470813 $T=277285 40770 1 0 $X=276885 $Y=39800
X794 22 VIA1_C_CDNS_7194277470813 $T=278825 38490 1 0 $X=278425 $Y=37520
X795 14 VIA1_C_CDNS_7194277470813 $T=280365 40770 1 0 $X=279965 $Y=39800
X796 22 VIA1_C_CDNS_7194277470813 $T=281905 38490 1 0 $X=281505 $Y=37520
X797 14 VIA1_C_CDNS_7194277470813 $T=283445 40770 1 0 $X=283045 $Y=39800
X798 22 VIA1_C_CDNS_7194277470813 $T=284985 38490 1 0 $X=284585 $Y=37520
X799 14 VIA1_C_CDNS_7194277470813 $T=286525 40770 1 0 $X=286125 $Y=39800
X800 22 VIA1_C_CDNS_7194277470813 $T=288065 38490 1 0 $X=287665 $Y=37520
X801 14 VIA1_C_CDNS_7194277470813 $T=289605 40770 1 0 $X=289205 $Y=39800
X802 22 VIA1_C_CDNS_7194277470813 $T=291145 38490 1 0 $X=290745 $Y=37520
X803 14 VIA1_C_CDNS_7194277470813 $T=292685 40770 1 0 $X=292285 $Y=39800
X804 22 VIA1_C_CDNS_7194277470813 $T=294225 38490 1 0 $X=293825 $Y=37520
X805 14 VIA1_C_CDNS_7194277470813 $T=295765 40770 1 0 $X=295365 $Y=39800
X806 15 VIA1_C_CDNS_7194277470813 $T=302300 40770 1 0 $X=301900 $Y=39800
X807 22 VIA1_C_CDNS_7194277470813 $T=303840 38490 1 0 $X=303440 $Y=37520
X808 15 VIA1_C_CDNS_7194277470813 $T=305380 40770 1 0 $X=304980 $Y=39800
X809 22 VIA1_C_CDNS_7194277470813 $T=306920 38490 1 0 $X=306520 $Y=37520
X810 15 VIA1_C_CDNS_7194277470813 $T=308460 40770 1 0 $X=308060 $Y=39800
X811 22 VIA1_C_CDNS_7194277470813 $T=310000 38490 1 0 $X=309600 $Y=37520
X812 15 VIA1_C_CDNS_7194277470813 $T=311540 40770 1 0 $X=311140 $Y=39800
X813 22 VIA1_C_CDNS_7194277470813 $T=313080 38490 1 0 $X=312680 $Y=37520
X814 15 VIA1_C_CDNS_7194277470813 $T=314620 40770 1 0 $X=314220 $Y=39800
X815 22 VIA1_C_CDNS_7194277470813 $T=316160 38490 1 0 $X=315760 $Y=37520
X816 15 VIA1_C_CDNS_7194277470813 $T=317700 40770 1 0 $X=317300 $Y=39800
X817 22 VIA1_C_CDNS_7194277470813 $T=319240 38490 1 0 $X=318840 $Y=37520
X818 15 VIA1_C_CDNS_7194277470813 $T=320780 40770 1 0 $X=320380 $Y=39800
X819 22 VIA1_C_CDNS_7194277470813 $T=322320 38490 1 0 $X=321920 $Y=37520
X820 15 VIA1_C_CDNS_7194277470813 $T=323860 40770 1 0 $X=323460 $Y=39800
X821 22 VIA1_C_CDNS_7194277470813 $T=325400 38490 1 0 $X=325000 $Y=37520
X822 15 VIA1_C_CDNS_7194277470813 $T=326940 40770 1 0 $X=326540 $Y=39800
X823 16 VIA1_C_CDNS_7194277470813 $T=333065 40770 1 0 $X=332665 $Y=39800
X824 22 VIA1_C_CDNS_7194277470813 $T=334605 38490 1 0 $X=334205 $Y=37520
X825 16 VIA1_C_CDNS_7194277470813 $T=336145 40770 1 0 $X=335745 $Y=39800
X826 22 VIA1_C_CDNS_7194277470813 $T=337685 38490 1 0 $X=337285 $Y=37520
X827 16 VIA1_C_CDNS_7194277470813 $T=339225 40770 1 0 $X=338825 $Y=39800
X828 22 VIA1_C_CDNS_7194277470813 $T=340765 38490 1 0 $X=340365 $Y=37520
X829 16 VIA1_C_CDNS_7194277470813 $T=342305 40770 1 0 $X=341905 $Y=39800
X830 22 VIA1_C_CDNS_7194277470813 $T=343845 38490 1 0 $X=343445 $Y=37520
X831 16 VIA1_C_CDNS_7194277470813 $T=345385 40770 1 0 $X=344985 $Y=39800
X832 20 VIA1_C_CDNS_7194277470813 $T=351530 40770 1 0 $X=351130 $Y=39800
X833 22 VIA1_C_CDNS_7194277470813 $T=353070 38490 1 0 $X=352670 $Y=37520
X834 20 VIA1_C_CDNS_7194277470813 $T=354610 40770 1 0 $X=354210 $Y=39800
X835 22 VIA1_C_CDNS_7194277470813 $T=356150 38490 1 0 $X=355750 $Y=37520
X836 20 VIA1_C_CDNS_7194277470813 $T=357690 40770 1 0 $X=357290 $Y=39800
X837 17 VIA1_C_CDNS_7194277470813 $T=363865 40770 1 0 $X=363465 $Y=39800
X838 22 VIA1_C_CDNS_7194277470813 $T=365405 38490 1 0 $X=365005 $Y=37520
X839 17 VIA1_C_CDNS_7194277470813 $T=366945 40770 1 0 $X=366545 $Y=39800
X840 19 VIA1_C_CDNS_7194277470813 $T=373240 40770 1 0 $X=372840 $Y=39800
X841 22 VIA1_C_CDNS_7194277470813 $T=374780 38490 1 0 $X=374380 $Y=37520
X842 4 VIA2_C_CDNS_7194277470814 $T=10890 144880 0 0 $X=10180 $Y=144220
X843 4 VIA2_C_CDNS_7194277470814 $T=10890 177040 0 0 $X=10180 $Y=176380
X844 10 VIA2_C_CDNS_7194277470814 $T=41770 143100 0 0 $X=41060 $Y=142440
X845 10 VIA2_C_CDNS_7194277470814 $T=41770 175260 0 0 $X=41060 $Y=174600
X846 5 VIA1_C_CDNS_7194277470816 $T=79820 146660 0 0 $X=78380 $Y=146470
X847 5 VIA1_C_CDNS_7194277470816 $T=79820 173480 0 0 $X=78380 $Y=173290
X848 5 VIA1_C_CDNS_7194277470816 $T=91060 146660 0 0 $X=89620 $Y=146470
X849 5 VIA1_C_CDNS_7194277470816 $T=91060 173480 0 0 $X=89620 $Y=173290
X850 5 VIA1_C_CDNS_7194277470816 $T=102300 146660 0 0 $X=100860 $Y=146470
X851 5 VIA1_C_CDNS_7194277470816 $T=102300 173480 0 0 $X=100860 $Y=173290
X852 5 VIA1_C_CDNS_7194277470816 $T=113540 146660 0 0 $X=112100 $Y=146470
X853 5 VIA1_C_CDNS_7194277470816 $T=113540 173480 0 0 $X=112100 $Y=173290
X854 5 VIA1_C_CDNS_7194277470816 $T=124780 146660 0 0 $X=123340 $Y=146470
X855 5 VIA1_C_CDNS_7194277470816 $T=124780 173480 0 0 $X=123340 $Y=173290
X856 5 VIA1_C_CDNS_7194277470816 $T=136020 146660 0 0 $X=134580 $Y=146470
X857 5 VIA1_C_CDNS_7194277470816 $T=136020 173480 0 0 $X=134580 $Y=173290
X858 5 VIA1_C_CDNS_7194277470816 $T=147260 146660 0 0 $X=145820 $Y=146470
X859 5 VIA1_C_CDNS_7194277470816 $T=147260 173480 0 0 $X=145820 $Y=173290
X860 5 VIA1_C_CDNS_7194277470816 $T=158500 146660 0 0 $X=157060 $Y=146470
X861 5 VIA1_C_CDNS_7194277470816 $T=158500 173480 0 0 $X=157060 $Y=173290
X862 13 VIA2_C_CDNS_7194277470817 $T=70100 98685 0 0 $X=69960 $Y=97975
X863 13 VIA2_C_CDNS_7194277470817 $T=70100 126585 0 0 $X=69960 $Y=125875
X864 13 VIA2_C_CDNS_7194277470817 $T=71370 98685 0 0 $X=71230 $Y=97975
X865 13 VIA2_C_CDNS_7194277470817 $T=71370 126585 0 0 $X=71230 $Y=125875
X866 13 VIA2_C_CDNS_7194277470817 $T=72640 98685 0 0 $X=72500 $Y=97975
X867 13 VIA2_C_CDNS_7194277470817 $T=72640 126585 0 0 $X=72500 $Y=125875
X868 13 VIA2_C_CDNS_7194277470817 $T=73500 98685 0 0 $X=73360 $Y=97975
X869 13 VIA2_C_CDNS_7194277470817 $T=73500 126585 0 0 $X=73360 $Y=125875
X870 13 VIA2_C_CDNS_7194277470817 $T=74770 98685 0 0 $X=74630 $Y=97975
X871 13 VIA2_C_CDNS_7194277470817 $T=74770 126585 0 0 $X=74630 $Y=125875
X872 6 VIA2_C_CDNS_7194277470817 $T=76040 96905 0 0 $X=75900 $Y=96195
X873 7 VIA2_C_CDNS_7194277470817 $T=76040 128365 0 0 $X=75900 $Y=127655
X874 13 VIA2_C_CDNS_7194277470817 $T=76900 98685 0 0 $X=76760 $Y=97975
X875 13 VIA2_C_CDNS_7194277470817 $T=76900 126585 0 0 $X=76760 $Y=125875
X876 13 VIA2_C_CDNS_7194277470817 $T=78170 98685 0 0 $X=78030 $Y=97975
X877 13 VIA2_C_CDNS_7194277470817 $T=78170 126585 0 0 $X=78030 $Y=125875
X878 7 VIA2_C_CDNS_7194277470817 $T=79440 95125 0 0 $X=79300 $Y=94415
X879 6 VIA2_C_CDNS_7194277470817 $T=79440 130145 0 0 $X=79300 $Y=129435
X880 13 VIA2_C_CDNS_7194277470817 $T=80300 98685 0 0 $X=80160 $Y=97975
X881 13 VIA2_C_CDNS_7194277470817 $T=80300 126585 0 0 $X=80160 $Y=125875
X882 13 VIA2_C_CDNS_7194277470817 $T=81570 98685 0 0 $X=81430 $Y=97975
X883 13 VIA2_C_CDNS_7194277470817 $T=81570 126585 0 0 $X=81430 $Y=125875
X884 6 VIA2_C_CDNS_7194277470817 $T=82840 96905 0 0 $X=82700 $Y=96195
X885 7 VIA2_C_CDNS_7194277470817 $T=82840 128365 0 0 $X=82700 $Y=127655
X886 13 VIA2_C_CDNS_7194277470817 $T=83700 98685 0 0 $X=83560 $Y=97975
X887 13 VIA2_C_CDNS_7194277470817 $T=83700 126585 0 0 $X=83560 $Y=125875
X888 13 VIA2_C_CDNS_7194277470817 $T=84970 98685 0 0 $X=84830 $Y=97975
X889 13 VIA2_C_CDNS_7194277470817 $T=84970 126585 0 0 $X=84830 $Y=125875
X890 7 VIA2_C_CDNS_7194277470817 $T=86240 95125 0 0 $X=86100 $Y=94415
X891 6 VIA2_C_CDNS_7194277470817 $T=86240 130145 0 0 $X=86100 $Y=129435
X892 13 VIA2_C_CDNS_7194277470817 $T=87100 98685 0 0 $X=86960 $Y=97975
X893 13 VIA2_C_CDNS_7194277470817 $T=87100 126585 0 0 $X=86960 $Y=125875
X894 13 VIA2_C_CDNS_7194277470817 $T=88370 98685 0 0 $X=88230 $Y=97975
X895 13 VIA2_C_CDNS_7194277470817 $T=88370 126585 0 0 $X=88230 $Y=125875
X896 6 VIA2_C_CDNS_7194277470817 $T=89640 96905 0 0 $X=89500 $Y=96195
X897 7 VIA2_C_CDNS_7194277470817 $T=89640 128365 0 0 $X=89500 $Y=127655
X898 13 VIA2_C_CDNS_7194277470817 $T=90500 98685 0 0 $X=90360 $Y=97975
X899 13 VIA2_C_CDNS_7194277470817 $T=90500 126585 0 0 $X=90360 $Y=125875
X900 13 VIA2_C_CDNS_7194277470817 $T=91770 98685 0 0 $X=91630 $Y=97975
X901 13 VIA2_C_CDNS_7194277470817 $T=91770 126585 0 0 $X=91630 $Y=125875
X902 7 VIA2_C_CDNS_7194277470817 $T=93040 95125 0 0 $X=92900 $Y=94415
X903 6 VIA2_C_CDNS_7194277470817 $T=93040 130145 0 0 $X=92900 $Y=129435
X904 13 VIA2_C_CDNS_7194277470817 $T=93900 98685 0 0 $X=93760 $Y=97975
X905 13 VIA2_C_CDNS_7194277470817 $T=93900 126585 0 0 $X=93760 $Y=125875
X906 13 VIA2_C_CDNS_7194277470817 $T=95170 98685 0 0 $X=95030 $Y=97975
X907 13 VIA2_C_CDNS_7194277470817 $T=95170 126585 0 0 $X=95030 $Y=125875
X908 6 VIA2_C_CDNS_7194277470817 $T=96440 96905 0 0 $X=96300 $Y=96195
X909 7 VIA2_C_CDNS_7194277470817 $T=96440 128365 0 0 $X=96300 $Y=127655
X910 13 VIA2_C_CDNS_7194277470817 $T=97300 98685 0 0 $X=97160 $Y=97975
X911 13 VIA2_C_CDNS_7194277470817 $T=97300 126585 0 0 $X=97160 $Y=125875
X912 13 VIA2_C_CDNS_7194277470817 $T=98570 98685 0 0 $X=98430 $Y=97975
X913 13 VIA2_C_CDNS_7194277470817 $T=98570 126585 0 0 $X=98430 $Y=125875
X914 7 VIA2_C_CDNS_7194277470817 $T=99840 95125 0 0 $X=99700 $Y=94415
X915 6 VIA2_C_CDNS_7194277470817 $T=99840 130145 0 0 $X=99700 $Y=129435
X916 13 VIA2_C_CDNS_7194277470817 $T=100700 98685 0 0 $X=100560 $Y=97975
X917 13 VIA2_C_CDNS_7194277470817 $T=100700 126585 0 0 $X=100560 $Y=125875
X918 13 VIA2_C_CDNS_7194277470817 $T=101970 98685 0 0 $X=101830 $Y=97975
X919 13 VIA2_C_CDNS_7194277470817 $T=101970 126585 0 0 $X=101830 $Y=125875
X920 6 VIA2_C_CDNS_7194277470817 $T=103240 96905 0 0 $X=103100 $Y=96195
X921 7 VIA2_C_CDNS_7194277470817 $T=103240 128365 0 0 $X=103100 $Y=127655
X922 13 VIA2_C_CDNS_7194277470817 $T=104100 98685 0 0 $X=103960 $Y=97975
X923 13 VIA2_C_CDNS_7194277470817 $T=104100 126585 0 0 $X=103960 $Y=125875
X924 13 VIA2_C_CDNS_7194277470817 $T=105370 98685 0 0 $X=105230 $Y=97975
X925 13 VIA2_C_CDNS_7194277470817 $T=105370 126585 0 0 $X=105230 $Y=125875
X926 7 VIA2_C_CDNS_7194277470817 $T=106640 95125 0 0 $X=106500 $Y=94415
X927 6 VIA2_C_CDNS_7194277470817 $T=106640 130145 0 0 $X=106500 $Y=129435
X928 13 VIA2_C_CDNS_7194277470817 $T=107500 98685 0 0 $X=107360 $Y=97975
X929 13 VIA2_C_CDNS_7194277470817 $T=107500 126585 0 0 $X=107360 $Y=125875
X930 13 VIA2_C_CDNS_7194277470817 $T=108770 98685 0 0 $X=108630 $Y=97975
X931 13 VIA2_C_CDNS_7194277470817 $T=108770 126585 0 0 $X=108630 $Y=125875
X932 6 VIA2_C_CDNS_7194277470817 $T=110040 96905 0 0 $X=109900 $Y=96195
X933 7 VIA2_C_CDNS_7194277470817 $T=110040 128365 0 0 $X=109900 $Y=127655
X934 13 VIA2_C_CDNS_7194277470817 $T=110900 98685 0 0 $X=110760 $Y=97975
X935 13 VIA2_C_CDNS_7194277470817 $T=110900 126585 0 0 $X=110760 $Y=125875
X936 13 VIA2_C_CDNS_7194277470817 $T=112170 98685 0 0 $X=112030 $Y=97975
X937 13 VIA2_C_CDNS_7194277470817 $T=112170 126585 0 0 $X=112030 $Y=125875
X938 7 VIA2_C_CDNS_7194277470817 $T=113440 95125 0 0 $X=113300 $Y=94415
X939 6 VIA2_C_CDNS_7194277470817 $T=113440 130145 0 0 $X=113300 $Y=129435
X940 13 VIA2_C_CDNS_7194277470817 $T=114300 98685 0 0 $X=114160 $Y=97975
X941 13 VIA2_C_CDNS_7194277470817 $T=114300 126585 0 0 $X=114160 $Y=125875
X942 13 VIA2_C_CDNS_7194277470817 $T=115570 98685 0 0 $X=115430 $Y=97975
X943 13 VIA2_C_CDNS_7194277470817 $T=115570 126585 0 0 $X=115430 $Y=125875
X944 6 VIA2_C_CDNS_7194277470817 $T=116840 96905 0 0 $X=116700 $Y=96195
X945 7 VIA2_C_CDNS_7194277470817 $T=116840 128365 0 0 $X=116700 $Y=127655
X946 13 VIA2_C_CDNS_7194277470817 $T=117700 98685 0 0 $X=117560 $Y=97975
X947 13 VIA2_C_CDNS_7194277470817 $T=117700 126585 0 0 $X=117560 $Y=125875
X948 13 VIA2_C_CDNS_7194277470817 $T=118970 98685 0 0 $X=118830 $Y=97975
X949 13 VIA2_C_CDNS_7194277470817 $T=118970 126585 0 0 $X=118830 $Y=125875
X950 7 VIA2_C_CDNS_7194277470817 $T=120240 95125 0 0 $X=120100 $Y=94415
X951 6 VIA2_C_CDNS_7194277470817 $T=120240 130145 0 0 $X=120100 $Y=129435
X952 13 VIA2_C_CDNS_7194277470817 $T=121100 98685 0 0 $X=120960 $Y=97975
X953 13 VIA2_C_CDNS_7194277470817 $T=121100 126585 0 0 $X=120960 $Y=125875
X954 13 VIA2_C_CDNS_7194277470817 $T=122370 98685 0 0 $X=122230 $Y=97975
X955 13 VIA2_C_CDNS_7194277470817 $T=122370 126585 0 0 $X=122230 $Y=125875
X956 6 VIA2_C_CDNS_7194277470817 $T=123640 96905 0 0 $X=123500 $Y=96195
X957 7 VIA2_C_CDNS_7194277470817 $T=123640 128365 0 0 $X=123500 $Y=127655
X958 13 VIA2_C_CDNS_7194277470817 $T=124500 98685 0 0 $X=124360 $Y=97975
X959 13 VIA2_C_CDNS_7194277470817 $T=124500 126585 0 0 $X=124360 $Y=125875
X960 13 VIA2_C_CDNS_7194277470817 $T=125770 98685 0 0 $X=125630 $Y=97975
X961 13 VIA2_C_CDNS_7194277470817 $T=125770 126585 0 0 $X=125630 $Y=125875
X962 7 VIA2_C_CDNS_7194277470817 $T=127040 95125 0 0 $X=126900 $Y=94415
X963 6 VIA2_C_CDNS_7194277470817 $T=127040 130145 0 0 $X=126900 $Y=129435
X964 13 VIA2_C_CDNS_7194277470817 $T=127900 98685 0 0 $X=127760 $Y=97975
X965 13 VIA2_C_CDNS_7194277470817 $T=127900 126585 0 0 $X=127760 $Y=125875
X966 13 VIA2_C_CDNS_7194277470817 $T=129170 98685 0 0 $X=129030 $Y=97975
X967 13 VIA2_C_CDNS_7194277470817 $T=129170 126585 0 0 $X=129030 $Y=125875
X968 13 VIA2_C_CDNS_7194277470817 $T=130440 98685 0 0 $X=130300 $Y=97975
X969 13 VIA2_C_CDNS_7194277470817 $T=130440 126585 0 0 $X=130300 $Y=125875
X970 13 VIA1_C_CDNS_7194277470818 $T=71370 100245 0 0 $X=70920 $Y=100105
X971 13 VIA1_C_CDNS_7194277470818 $T=71370 125025 0 0 $X=70920 $Y=124885
X972 13 VIA1_C_CDNS_7194277470818 $T=74770 100245 0 0 $X=74320 $Y=100105
X973 13 VIA1_C_CDNS_7194277470818 $T=74770 125025 0 0 $X=74320 $Y=124885
X974 13 VIA1_C_CDNS_7194277470818 $T=78170 100245 0 0 $X=77720 $Y=100105
X975 13 VIA1_C_CDNS_7194277470818 $T=78170 125025 0 0 $X=77720 $Y=124885
X976 13 VIA1_C_CDNS_7194277470818 $T=81570 100245 0 0 $X=81120 $Y=100105
X977 13 VIA1_C_CDNS_7194277470818 $T=81570 125025 0 0 $X=81120 $Y=124885
X978 13 VIA1_C_CDNS_7194277470818 $T=84970 100245 0 0 $X=84520 $Y=100105
X979 13 VIA1_C_CDNS_7194277470818 $T=84970 125025 0 0 $X=84520 $Y=124885
X980 13 VIA1_C_CDNS_7194277470818 $T=88370 100245 0 0 $X=87920 $Y=100105
X981 13 VIA1_C_CDNS_7194277470818 $T=88370 125025 0 0 $X=87920 $Y=124885
X982 13 VIA1_C_CDNS_7194277470818 $T=91770 100245 0 0 $X=91320 $Y=100105
X983 13 VIA1_C_CDNS_7194277470818 $T=91770 125025 0 0 $X=91320 $Y=124885
X984 13 VIA1_C_CDNS_7194277470818 $T=95170 100245 0 0 $X=94720 $Y=100105
X985 13 VIA1_C_CDNS_7194277470818 $T=95170 125025 0 0 $X=94720 $Y=124885
X986 13 VIA1_C_CDNS_7194277470818 $T=98570 100245 0 0 $X=98120 $Y=100105
X987 13 VIA1_C_CDNS_7194277470818 $T=98570 125025 0 0 $X=98120 $Y=124885
X988 13 VIA1_C_CDNS_7194277470818 $T=101970 100245 0 0 $X=101520 $Y=100105
X989 13 VIA1_C_CDNS_7194277470818 $T=101970 125025 0 0 $X=101520 $Y=124885
X990 13 VIA1_C_CDNS_7194277470818 $T=105370 100245 0 0 $X=104920 $Y=100105
X991 13 VIA1_C_CDNS_7194277470818 $T=105370 125025 0 0 $X=104920 $Y=124885
X992 13 VIA1_C_CDNS_7194277470818 $T=108770 100245 0 0 $X=108320 $Y=100105
X993 13 VIA1_C_CDNS_7194277470818 $T=108770 125025 0 0 $X=108320 $Y=124885
X994 13 VIA1_C_CDNS_7194277470818 $T=112170 100245 0 0 $X=111720 $Y=100105
X995 13 VIA1_C_CDNS_7194277470818 $T=112170 125025 0 0 $X=111720 $Y=124885
X996 13 VIA1_C_CDNS_7194277470818 $T=115570 100245 0 0 $X=115120 $Y=100105
X997 13 VIA1_C_CDNS_7194277470818 $T=115570 125025 0 0 $X=115120 $Y=124885
X998 13 VIA1_C_CDNS_7194277470818 $T=118970 100245 0 0 $X=118520 $Y=100105
X999 13 VIA1_C_CDNS_7194277470818 $T=118970 125025 0 0 $X=118520 $Y=124885
X1000 13 VIA1_C_CDNS_7194277470818 $T=122370 100245 0 0 $X=121920 $Y=100105
X1001 13 VIA1_C_CDNS_7194277470818 $T=122370 125025 0 0 $X=121920 $Y=124885
X1002 13 VIA1_C_CDNS_7194277470818 $T=125770 100245 0 0 $X=125320 $Y=100105
X1003 13 VIA1_C_CDNS_7194277470818 $T=125770 125025 0 0 $X=125320 $Y=124885
X1004 13 VIA1_C_CDNS_7194277470818 $T=129170 100245 0 0 $X=128720 $Y=100105
X1005 13 VIA1_C_CDNS_7194277470818 $T=129170 125025 0 0 $X=128720 $Y=124885
X1006 7 VIA3_C_CDNS_7194277470819 $T=63650 95125 0 0 $X=62680 $Y=94465
X1007 7 VIA3_C_CDNS_7194277470819 $T=63650 128365 0 0 $X=62680 $Y=127705
X1008 6 VIA3_C_CDNS_7194277470819 $T=65930 96905 0 0 $X=64960 $Y=96245
X1009 6 VIA3_C_CDNS_7194277470819 $T=65930 130145 0 0 $X=64960 $Y=129485
X1010 13 VIA3_C_CDNS_7194277470819 $T=68210 98685 0 0 $X=67240 $Y=98025
X1011 13 VIA3_C_CDNS_7194277470819 $T=68210 126585 0 0 $X=67240 $Y=125925
X1012 13 VIA3_C_CDNS_7194277470819 $T=132330 98685 0 0 $X=131360 $Y=98025
X1013 13 VIA3_C_CDNS_7194277470819 $T=132330 126585 0 0 $X=131360 $Y=125925
X1014 7 VIA3_C_CDNS_7194277470819 $T=134610 95125 0 0 $X=133640 $Y=94465
X1015 7 VIA3_C_CDNS_7194277470819 $T=134610 128365 0 0 $X=133640 $Y=127705
X1016 6 VIA3_C_CDNS_7194277470819 $T=136890 96905 0 0 $X=135920 $Y=96245
X1017 6 VIA3_C_CDNS_7194277470819 $T=136890 130145 0 0 $X=135920 $Y=129485
X1018 23 VIA2_C_CDNS_7194277470820 $T=74460 112235 0 0 $X=74320 $Y=112045
X1019 21 VIA2_C_CDNS_7194277470820 $T=75080 113015 0 0 $X=74940 $Y=112825
X1020 23 VIA2_C_CDNS_7194277470820 $T=78170 112235 0 0 $X=78030 $Y=112045
X1021 21 VIA2_C_CDNS_7194277470820 $T=78170 113015 0 0 $X=78030 $Y=112825
X1022 23 VIA2_C_CDNS_7194277470820 $T=81260 112235 0 0 $X=81120 $Y=112045
X1023 21 VIA2_C_CDNS_7194277470820 $T=81880 113015 0 0 $X=81740 $Y=112825
X1024 23 VIA2_C_CDNS_7194277470820 $T=84970 112235 0 0 $X=84830 $Y=112045
X1025 21 VIA2_C_CDNS_7194277470820 $T=84970 113015 0 0 $X=84830 $Y=112825
X1026 23 VIA2_C_CDNS_7194277470820 $T=88060 112235 0 0 $X=87920 $Y=112045
X1027 21 VIA2_C_CDNS_7194277470820 $T=88680 113015 0 0 $X=88540 $Y=112825
X1028 23 VIA2_C_CDNS_7194277470820 $T=91770 112235 0 0 $X=91630 $Y=112045
X1029 21 VIA2_C_CDNS_7194277470820 $T=91770 113015 0 0 $X=91630 $Y=112825
X1030 23 VIA2_C_CDNS_7194277470820 $T=94860 112235 0 0 $X=94720 $Y=112045
X1031 21 VIA2_C_CDNS_7194277470820 $T=95480 113015 0 0 $X=95340 $Y=112825
X1032 23 VIA2_C_CDNS_7194277470820 $T=98570 112235 0 0 $X=98430 $Y=112045
X1033 21 VIA2_C_CDNS_7194277470820 $T=98570 113015 0 0 $X=98430 $Y=112825
X1034 23 VIA2_C_CDNS_7194277470820 $T=101660 112235 0 0 $X=101520 $Y=112045
X1035 21 VIA2_C_CDNS_7194277470820 $T=102280 113015 0 0 $X=102140 $Y=112825
X1036 23 VIA2_C_CDNS_7194277470820 $T=105370 112235 0 0 $X=105230 $Y=112045
X1037 21 VIA2_C_CDNS_7194277470820 $T=105370 113015 0 0 $X=105230 $Y=112825
X1038 23 VIA2_C_CDNS_7194277470820 $T=108460 112235 0 0 $X=108320 $Y=112045
X1039 21 VIA2_C_CDNS_7194277470820 $T=109080 113015 0 0 $X=108940 $Y=112825
X1040 23 VIA2_C_CDNS_7194277470820 $T=112170 112235 0 0 $X=112030 $Y=112045
X1041 21 VIA2_C_CDNS_7194277470820 $T=112170 113015 0 0 $X=112030 $Y=112825
X1042 23 VIA2_C_CDNS_7194277470820 $T=115260 112235 0 0 $X=115120 $Y=112045
X1043 21 VIA2_C_CDNS_7194277470820 $T=115880 113015 0 0 $X=115740 $Y=112825
X1044 23 VIA2_C_CDNS_7194277470820 $T=118970 112235 0 0 $X=118830 $Y=112045
X1045 21 VIA2_C_CDNS_7194277470820 $T=118970 113015 0 0 $X=118830 $Y=112825
X1046 23 VIA2_C_CDNS_7194277470820 $T=122060 112235 0 0 $X=121920 $Y=112045
X1047 21 VIA2_C_CDNS_7194277470820 $T=122680 113015 0 0 $X=122540 $Y=112825
X1048 23 VIA2_C_CDNS_7194277470820 $T=125770 112235 0 0 $X=125630 $Y=112045
X1049 21 VIA2_C_CDNS_7194277470820 $T=125770 113015 0 0 $X=125630 $Y=112825
X1050 24 VIA1_C_CDNS_7194277470822 $T=89720 58980 0 0 $X=88970 $Y=58750
X1051 24 VIA1_C_CDNS_7194277470822 $T=89825 61565 0 90 $X=89595 $Y=60815
X1052 5 VIA1_C_CDNS_7194277470823 $T=90930 69330 0 0 $X=88880 $Y=68840
X1053 5 VIA1_C_CDNS_7194277470823 $T=90930 73450 0 0 $X=88880 $Y=72960
X1054 11 VIA1_C_CDNS_7194277470824 $T=300690 18770 0 0 $X=299160 $Y=17760
X1055 11 VIA1_C_CDNS_7194277470824 $T=306120 19025 0 0 $X=304590 $Y=18015
X1056 2 VIA2_C_CDNS_7194277470825 $T=7140 58145 0 0 $X=5610 $Y=57395
X1057 1 VIA2_C_CDNS_7194277470825 $T=17075 56365 0 0 $X=15545 $Y=55615
X1058 5 11 VIA1_C_CDNS_7194277470826 $T=13915 179845 0 0 $X=8745 $Y=178835
X1059 5 11 VIA1_C_CDNS_7194277470826 $T=38730 179845 0 0 $X=33560 $Y=178835
X1060 5 11 VIA1_C_CDNS_7194277470826 $T=54060 179845 0 0 $X=48890 $Y=178835
X1061 5 11 VIA1_C_CDNS_7194277470826 $T=169780 179845 0 0 $X=164610 $Y=178835
X1062 5 11 VIA1_C_CDNS_7194277470826 $T=202645 179775 0 0 $X=197475 $Y=178765
X1063 5 11 VIA1_C_CDNS_7194277470826 $T=375600 179775 0 0 $X=370430 $Y=178765
X1064 5 11 VIA2_C_CDNS_7194277470827 $T=202645 179775 0 0 $X=197475 $Y=178765
X1065 5 11 VIA2_C_CDNS_7194277470827 $T=375600 179775 0 0 $X=370430 $Y=178765
X1066 5 VIA1_C_CDNS_7194277470828 $T=57370 119810 0 0 $X=56880 $Y=116720
X1067 5 VIA1_C_CDNS_7194277470828 $T=67590 119810 0 0 $X=67100 $Y=116720
X1068 5 VIA1_C_CDNS_7194277470828 $T=132950 119810 0 0 $X=132460 $Y=116720
X1069 5 VIA1_C_CDNS_7194277470828 $T=143170 119810 0 0 $X=142680 $Y=116720
X1070 21 VIA1_C_CDNS_7194277470832 $T=75215 41040 0 0 $X=74725 $Y=38990
X1071 22 VIA1_C_CDNS_7194277470832 $T=185295 41010 0 0 $X=184805 $Y=38960
X1072 18 VIA2_C_CDNS_7194277470833 $T=225125 38490 0 0 $X=224125 $Y=37490
X1073 14 VIA2_C_CDNS_7194277470833 $T=305715 12525 0 0 $X=304715 $Y=11525
X1074 15 VIA2_C_CDNS_7194277470833 $T=318935 12525 0 0 $X=317935 $Y=11525
X1075 16 VIA2_C_CDNS_7194277470833 $T=328195 12525 0 0 $X=327195 $Y=11525
X1076 20 VIA2_C_CDNS_7194277470833 $T=337455 12525 0 0 $X=336455 $Y=11525
X1077 17 VIA2_C_CDNS_7194277470833 $T=346715 12525 0 0 $X=345715 $Y=11525
X1078 19 VIA2_C_CDNS_7194277470833 $T=355975 12525 0 0 $X=354975 $Y=11525
X1079 12 VIA2_C_CDNS_7194277470834 $T=63460 55465 0 0 $X=61410 $Y=54455
X1080 22 VIA2_C_CDNS_7194277470834 $T=247295 38480 0 0 $X=245245 $Y=37470
X1081 14 VIA2_C_CDNS_7194277470834 $T=294955 40780 0 0 $X=292905 $Y=39770
X1082 15 VIA2_C_CDNS_7194277470834 $T=303110 40780 0 0 $X=301060 $Y=39770
X1083 16 VIA2_C_CDNS_7194277470834 $T=344575 40780 0 0 $X=342525 $Y=39770
X1084 20 VIA2_C_CDNS_7194277470834 $T=356880 40780 0 0 $X=354830 $Y=39770
X1085 17 VIA2_C_CDNS_7194277470834 $T=365495 40780 0 0 $X=363445 $Y=39770
X1086 19 VIA2_C_CDNS_7194277470834 $T=374005 40780 0 0 $X=371955 $Y=39770
X1087 15 VIA3_C_CDNS_7194277470838 $T=303110 40780 0 0 $X=301060 $Y=39770
X1088 16 VIA3_C_CDNS_7194277470838 $T=344575 40780 0 0 $X=342525 $Y=39770
X1089 19 VIA3_C_CDNS_7194277470838 $T=374005 40780 0 0 $X=371955 $Y=39770
X1090 15 VIA3_C_CDNS_7194277470840 $T=195805 49055 0 0 $X=194805 $Y=48055
X1091 19 VIA3_C_CDNS_7194277470840 $T=377865 50400 0 0 $X=376865 $Y=49400
X1092 16 VIA3_C_CDNS_7194277470840 $T=386985 47530 0 0 $X=385985 $Y=46530
X1093 8 VIA1_C_CDNS_7194277470843 $T=151480 80915 0 0 $X=150730 $Y=78865
X1094 10 VIA1_C_CDNS_7194277470843 $T=151480 122460 0 0 $X=150730 $Y=120410
X1095 24 VIA2_C_CDNS_7194277470846 $T=89070 58460 0 0 $X=88320 $Y=57710
X1096 25 VIA2_C_CDNS_7194277470846 $T=307715 6345 0 0 $X=306965 $Y=5595
X1097 26 VIA2_C_CDNS_7194277470846 $T=316955 6345 0 0 $X=316205 $Y=5595
X1098 27 VIA2_C_CDNS_7194277470846 $T=326225 6345 0 0 $X=325475 $Y=5595
X1099 28 VIA2_C_CDNS_7194277470846 $T=335490 6345 0 0 $X=334740 $Y=5595
X1100 29 VIA2_C_CDNS_7194277470846 $T=344750 6345 0 0 $X=344000 $Y=5595
X1101 30 VIA2_C_CDNS_7194277470846 $T=354005 6345 0 0 $X=353255 $Y=5595
X1102 5 4 4 11 pe3_CDNS_719427747080 $T=15710 148580 0 0 $X=14200 $Y=147550
X1103 5 4 10 11 pe3_CDNS_719427747080 $T=26950 148580 0 0 $X=25440 $Y=147550
X1104 5 5 5 11 pe3_CDNS_719427747080 $T=56340 148580 0 0 $X=54830 $Y=147550
X1105 5 6 6 11 pe3_CDNS_719427747080 $T=67580 148580 0 0 $X=66070 $Y=147550
X1106 5 6 7 11 pe3_CDNS_719427747080 $T=78820 148580 0 0 $X=77310 $Y=147550
X1107 5 6 6 11 pe3_CDNS_719427747080 $T=90060 148580 0 0 $X=88550 $Y=147550
X1108 5 6 7 11 pe3_CDNS_719427747080 $T=101300 148580 0 0 $X=99790 $Y=147550
X1109 5 6 6 11 pe3_CDNS_719427747080 $T=112540 148580 0 0 $X=111030 $Y=147550
X1110 5 6 7 11 pe3_CDNS_719427747080 $T=123780 148580 0 0 $X=122270 $Y=147550
X1111 5 6 6 11 pe3_CDNS_719427747080 $T=135020 148580 0 0 $X=133510 $Y=147550
X1112 5 6 7 11 pe3_CDNS_719427747080 $T=146260 148580 0 0 $X=144750 $Y=147550
X1113 5 5 5 11 pe3_CDNS_719427747080 $T=157500 148580 0 0 $X=155990 $Y=147550
X1114 5 5 5 11 pe3_CDNS_719427747080 $T=362795 71115 1 0 $X=361285 $Y=60085
X1115 5 5 5 11 pe3_CDNS_719427747080 $T=362795 89915 1 0 $X=361285 $Y=78885
X1116 5 5 5 11 pe3_CDNS_719427747080 $T=362795 108715 1 0 $X=361285 $Y=97685
X1117 5 5 5 11 pe3_CDNS_719427747080 $T=362795 127515 1 0 $X=361285 $Y=116485
X1118 5 5 5 11 pe3_CDNS_719427747080 $T=362795 146315 1 0 $X=361285 $Y=135285
X1119 5 5 5 11 pe3_CDNS_719427747080 $T=362795 165115 1 0 $X=361285 $Y=154085
X1120 19 9 22 5 11 pe3_CDNS_719427747081 $T=373510 36320 1 0 $X=372000 $Y=25290
X1121 17 9 22 5 11 pe3_CDNS_719427747082 $T=364135 36320 1 0 $X=362625 $Y=25290
X1122 20 9 22 5 11 pe3_CDNS_719427747083 $T=351800 36320 1 0 $X=350290 $Y=25290
X1123 16 9 22 5 11 pe3_CDNS_719427747084 $T=333335 36320 1 0 $X=331825 $Y=25290
X1124 15 9 22 5 11 pe3_CDNS_719427747085 $T=302570 36320 1 0 $X=301060 $Y=25290
X1125 14 9 22 5 11 pe3_CDNS_719427747086 $T=246755 36320 1 0 $X=245245 $Y=25290
X1126 22 11 rpp1k1_3_CDNS_719427747087 $T=190390 9160 0 0 $X=185230 $Y=8940
X1127 18 9 21 5 11 pe3_CDNS_719427747088 $T=223935 36320 1 0 $X=222425 $Y=25290
X1128 21 11 rpp1k1_3_CDNS_719427747089 $T=80195 9200 0 0 $X=75035 $Y=8980
X1129 8 11 11 pe3_CDNS_7194277470810 $T=154675 76695 0 0 $X=153165 $Y=75665
X1130 9 8 11 pe3_CDNS_7194277470810 $T=154675 98175 0 0 $X=153165 $Y=97145
X1131 10 9 11 pe3_CDNS_7194277470810 $T=154675 119125 0 0 $X=153165 $Y=118095
X1132 5 24 31 11 pe3_CDNS_7194277470811 $T=91085 67915 1 0 $X=90175 $Y=61345
X1133 14 25 11 5 pe3_CDNS_7194277470812 $T=307075 17335 1 0 $X=305565 $Y=6305
X1134 15 26 11 5 pe3_CDNS_7194277470812 $T=316335 17335 1 0 $X=314825 $Y=6305
X1135 16 27 11 5 pe3_CDNS_7194277470812 $T=325595 17335 1 0 $X=324085 $Y=6305
X1136 20 28 11 5 pe3_CDNS_7194277470812 $T=334855 17335 1 0 $X=333345 $Y=6305
X1137 17 29 11 5 pe3_CDNS_7194277470812 $T=344115 17335 1 0 $X=342605 $Y=6305
X1138 19 30 11 5 pe3_CDNS_7194277470812 $T=353375 17335 1 0 $X=351865 $Y=6305
X1139 1 2 2 11 ne3_CDNS_7194277470813 $T=7715 59435 0 0 $X=6915 $Y=59035
X1140 3 2 4 11 ne3_CDNS_7194277470813 $T=34470 59435 0 0 $X=33670 $Y=59035
X1141 12 2 13 11 ne3_CDNS_7194277470813 $T=62205 59435 0 0 $X=61405 $Y=59035
X1142 11 11 11 ne3_CDNS_7194277470815 $T=11530 16320 0 0 $X=10730 $Y=15920
X1143 11 11 11 ne3_CDNS_7194277470815 $T=11530 38460 1 0 $X=10730 $Y=27890
X1144 11 1 12 ne3_CDNS_7194277470815 $T=14770 16320 0 0 $X=13970 $Y=15920
X1145 11 1 1 ne3_CDNS_7194277470815 $T=14770 38460 1 0 $X=13970 $Y=27890
X1146 11 1 3 ne3_CDNS_7194277470815 $T=18010 16320 0 0 $X=17210 $Y=15920
X1147 11 1 12 ne3_CDNS_7194277470815 $T=18010 38460 1 0 $X=17210 $Y=27890
X1148 11 1 1 ne3_CDNS_7194277470815 $T=21250 16320 0 0 $X=20450 $Y=15920
X1149 11 1 3 ne3_CDNS_7194277470815 $T=21250 38460 1 0 $X=20450 $Y=27890
X1150 11 1 12 ne3_CDNS_7194277470815 $T=24490 16320 0 0 $X=23690 $Y=15920
X1151 11 1 1 ne3_CDNS_7194277470815 $T=24490 38460 1 0 $X=23690 $Y=27890
X1152 11 1 3 ne3_CDNS_7194277470815 $T=27730 16320 0 0 $X=26930 $Y=15920
X1153 11 1 12 ne3_CDNS_7194277470815 $T=27730 38460 1 0 $X=26930 $Y=27890
X1154 11 1 1 ne3_CDNS_7194277470815 $T=30970 16320 0 0 $X=30170 $Y=15920
X1155 11 1 3 ne3_CDNS_7194277470815 $T=30970 38460 1 0 $X=30170 $Y=27890
X1156 11 1 12 ne3_CDNS_7194277470815 $T=34210 16320 0 0 $X=33410 $Y=15920
X1157 11 1 1 ne3_CDNS_7194277470815 $T=34210 38460 1 0 $X=33410 $Y=27890
X1158 11 1 3 ne3_CDNS_7194277470815 $T=37450 16320 0 0 $X=36650 $Y=15920
X1159 11 1 12 ne3_CDNS_7194277470815 $T=37450 38460 1 0 $X=36650 $Y=27890
X1160 11 1 1 ne3_CDNS_7194277470815 $T=40690 16320 0 0 $X=39890 $Y=15920
X1161 11 1 3 ne3_CDNS_7194277470815 $T=40690 38460 1 0 $X=39890 $Y=27890
X1162 11 1 12 ne3_CDNS_7194277470815 $T=43930 16320 0 0 $X=43130 $Y=15920
X1163 11 1 1 ne3_CDNS_7194277470815 $T=43930 38460 1 0 $X=43130 $Y=27890
X1164 11 1 3 ne3_CDNS_7194277470815 $T=47170 16320 0 0 $X=46370 $Y=15920
X1165 11 1 12 ne3_CDNS_7194277470815 $T=47170 38460 1 0 $X=46370 $Y=27890
X1166 11 1 1 ne3_CDNS_7194277470815 $T=50410 16320 0 0 $X=49610 $Y=15920
X1167 11 1 3 ne3_CDNS_7194277470815 $T=50410 38460 1 0 $X=49610 $Y=27890
X1168 11 11 11 ne3_CDNS_7194277470815 $T=53650 16320 0 0 $X=52850 $Y=15920
X1169 11 11 11 ne3_CDNS_7194277470815 $T=53650 38460 1 0 $X=52850 $Y=27890
X1170 5 11 pe3_CDNS_7194277470816 $T=362795 52315 1 0 $X=361285 $Y=49285
X1171 5 11 pe3_CDNS_7194277470816 $T=362795 175915 1 0 $X=361285 $Y=172885
X1172 11 31 1 ne3_CDNS_7194277470817 $T=96785 56345 0 0 $X=95985 $Y=55765
X1173 11 31 22 ne3_CDNS_7194277470817 $T=102390 56345 0 0 $X=101590 $Y=55765
X1174 11 24 31 ne3_CDNS_7194277470818 $T=91035 56560 0 0 $X=90235 $Y=56160
X1175 5 11 MASCO__A1 $T=203925 49285 0 0 $X=203925 $Y=49285
X1176 5 11 MASCO__A1 $T=203925 172885 0 0 $X=203925 $Y=172885
X1177 5 11 MASCO__A1 $T=226405 49285 0 0 $X=226405 $Y=49285
X1178 5 11 MASCO__A1 $T=226405 172885 0 0 $X=226405 $Y=172885
X1179 5 11 MASCO__A1 $T=248885 49285 0 0 $X=248885 $Y=49285
X1180 5 11 MASCO__A1 $T=248885 172885 0 0 $X=248885 $Y=172885
X1181 5 11 MASCO__A1 $T=271365 49285 0 0 $X=271365 $Y=49285
X1182 5 11 MASCO__A1 $T=271365 172885 0 0 $X=271365 $Y=172885
X1183 5 11 MASCO__A1 $T=293845 49285 0 0 $X=293845 $Y=49285
X1184 5 11 MASCO__A1 $T=293845 172885 0 0 $X=293845 $Y=172885
X1185 5 11 MASCO__A1 $T=316325 49285 0 0 $X=316325 $Y=49285
X1186 5 11 MASCO__A1 $T=316325 172885 0 0 $X=316325 $Y=172885
X1187 5 11 MASCO__A1 $T=338805 49285 0 0 $X=338805 $Y=49285
X1188 5 11 MASCO__A1 $T=338805 172885 0 0 $X=338805 $Y=172885
X1189 5 10 4 4 4 11 MASCO__A2 $T=14200 160530 0 0 $X=14200 $Y=160530
X1190 5 6 5 6 5 11 MASCO__A2 $T=144750 160530 0 0 $X=144750 $Y=160530
X1191 5 5 5 5 5 11 MASCO__A2 $T=338805 60085 0 0 $X=338805 $Y=60085
X1192 5 14 14 7 7 11 MASCO__A2 $T=338805 78885 0 0 $X=338805 $Y=78885
X1193 5 14 14 7 7 11 MASCO__A2 $T=338805 97685 0 0 $X=338805 $Y=97685
X1194 5 14 14 7 7 11 MASCO__A2 $T=338805 116485 0 0 $X=338805 $Y=116485
X1195 5 14 14 7 7 11 MASCO__A2 $T=338805 135285 0 0 $X=338805 $Y=135285
X1196 5 14 14 7 7 11 MASCO__A2 $T=338805 154085 0 0 $X=338805 $Y=154085
X1197 13 5 13 13 7 6 21 13 23 13
+ 11 MASCO__B5 $T=66310 96535 0 0 $X=66310 $Y=96535
X1198 13 5 6 7 7 6 21 23 23 21
+ 11 MASCO__B5 $T=73110 96535 0 0 $X=73110 $Y=96535
X1199 13 5 6 7 7 6 21 23 23 21
+ 11 MASCO__B5 $T=79910 96535 0 0 $X=79910 $Y=96535
X1200 13 5 6 7 7 6 21 23 23 21
+ 11 MASCO__B5 $T=86710 96535 0 0 $X=86710 $Y=96535
X1201 13 5 6 7 7 6 21 23 23 21
+ 11 MASCO__B5 $T=93510 96535 0 0 $X=93510 $Y=96535
X1202 13 5 6 7 7 6 21 23 23 21
+ 11 MASCO__B5 $T=100310 96535 0 0 $X=100310 $Y=96535
X1203 13 5 6 7 7 6 21 23 23 21
+ 11 MASCO__B5 $T=107110 96535 0 0 $X=107110 $Y=96535
X1204 13 5 6 7 7 6 21 23 23 21
+ 11 MASCO__B5 $T=113910 96535 0 0 $X=113910 $Y=96535
X1205 13 5 6 7 13 13 13 23 13 21
+ 11 MASCO__B5 $T=120710 96535 0 0 $X=120710 $Y=96535
X1206 5 5 6 7 6 7 5 11 MASCO__A6 $T=54830 160530 0 0 $X=54830 $Y=160530
X1207 5 6 6 7 6 7 6 11 MASCO__A6 $T=99790 160530 0 0 $X=99790 $Y=160530
X1208 5 5 7 14 15 15 5 11 MASCO__A6 $T=203925 60085 0 0 $X=203925 $Y=60085
X1209 5 5 7 14 15 16 5 11 MASCO__A6 $T=203925 78885 0 0 $X=203925 $Y=78885
X1210 5 5 7 14 15 16 5 11 MASCO__A6 $T=203925 97685 0 0 $X=203925 $Y=97685
X1211 5 5 7 14 15 16 5 11 MASCO__A6 $T=203925 116485 0 0 $X=203925 $Y=116485
X1212 5 5 7 14 15 16 5 11 MASCO__A6 $T=203925 135285 0 0 $X=203925 $Y=135285
X1213 5 5 7 14 14 14 5 11 MASCO__A6 $T=203925 154085 0 0 $X=203925 $Y=154085
X1214 5 15 7 15 18 14 7 11 MASCO__A6 $T=248885 60085 0 0 $X=248885 $Y=60085
X1215 5 18 7 20 20 18 7 11 MASCO__A6 $T=248885 78885 0 0 $X=248885 $Y=78885
X1216 5 17 7 18 19 18 7 11 MASCO__A6 $T=248885 97685 0 0 $X=248885 $Y=97685
X1217 5 18 7 17 18 16 7 11 MASCO__A6 $T=248885 116485 0 0 $X=248885 $Y=116485
X1218 5 18 7 20 20 18 7 11 MASCO__A6 $T=248885 135285 0 0 $X=248885 $Y=135285
X1219 5 14 7 14 15 15 7 11 MASCO__A6 $T=248885 154085 0 0 $X=248885 $Y=154085
X1220 5 14 5 5 5 5 7 11 MASCO__A6 $T=293845 60085 0 0 $X=293845 $Y=60085
X1221 5 16 7 15 14 14 7 11 MASCO__A6 $T=293845 78885 0 0 $X=293845 $Y=78885
X1222 5 16 7 15 14 14 7 11 MASCO__A6 $T=293845 97685 0 0 $X=293845 $Y=97685
X1223 5 15 7 15 14 14 7 11 MASCO__A6 $T=293845 116485 0 0 $X=293845 $Y=116485
X1224 5 16 7 15 14 14 7 11 MASCO__A6 $T=293845 135285 0 0 $X=293845 $Y=135285
X1225 5 15 7 18 14 14 7 11 MASCO__A6 $T=293845 154085 0 0 $X=293845 $Y=154085
D0 11 5 p_dnw AREA=7.95604e-10 PJ=0.00014876 perimeter=0.00014876 $X=8500 $Y=140710 $dt=3
D1 11 5 p_dnw AREA=2.14716e-09 PJ=0.0003306 perimeter=0.0003306 $X=48630 $Y=140710 $dt=3
D2 11 5 p_dnw AREA=3.11448e-11 PJ=3.188e-05 perimeter=3.188e-05 $X=88435 $Y=59745 $dt=3
D3 11 8 p_dnw AREA=1.97548e-10 PJ=8.944e-05 perimeter=8.944e-05 $X=151005 $Y=72505 $dt=3
D4 11 9 p_dnw AREA=1.97548e-10 PJ=8.944e-05 perimeter=8.944e-05 $X=151005 $Y=93985 $dt=3
D5 11 10 p_dnw AREA=1.97548e-10 PJ=8.944e-05 perimeter=8.944e-05 $X=151005 $Y=114935 $dt=3
D6 11 5 p_dnw AREA=1.47356e-08 PJ=0.0006944 perimeter=0.0006944 $X=181765 $Y=46865 $dt=3
D7 11 5 p_dnw AREA=1.65707e-09 PJ=0.00035483 perimeter=0.00035483 $X=220785 $Y=22870 $dt=3
D8 11 5 p_dnw AREA=6.02548e-10 PJ=0.00014223 perimeter=0.00014223 $X=303405 $Y=4665 $dt=3
D9 11 5 p_ddnw AREA=1.72778e-09 PJ=0.0002104 perimeter=0.0002104 $X=65040 $Y=95265 $dt=4
D10 13 5 p_dipdnwmv AREA=9.7703e-10 PJ=0.0001796 perimeter=0.0001796 $X=68890 $Y=99115 $dt=5
D11 11 5 p_dnw3 AREA=2.92576e-10 PJ=0 perimeter=0 $X=14200 $Y=147550 $dt=6
D12 11 5 p_dnw3 AREA=2.92576e-10 PJ=0 perimeter=0 $X=14200 $Y=160530 $dt=6
D13 11 5 p_dnw3 AREA=1.37701e-09 PJ=0 perimeter=0 $X=54830 $Y=147550 $dt=6
D14 11 5 p_dnw3 AREA=1.37701e-09 PJ=0 perimeter=0 $X=54830 $Y=160530 $dt=6
D15 11 5 p_dnw3 AREA=2.67592e-11 PJ=0 perimeter=0 $X=89575 $Y=60885 $dt=6
D16 11 5 p_dnw3 AREA=6.91743e-10 PJ=0 perimeter=0 $X=203925 $Y=49285 $dt=6
D17 11 5 p_dnw3 AREA=2.05478e-09 PJ=0 perimeter=0 $X=203925 $Y=60085 $dt=6
D18 11 5 p_dnw3 AREA=2.05478e-09 PJ=0 perimeter=0 $X=203925 $Y=78885 $dt=6
D19 11 5 p_dnw3 AREA=2.05478e-09 PJ=0 perimeter=0 $X=203925 $Y=97685 $dt=6
D20 11 5 p_dnw3 AREA=2.05478e-09 PJ=0 perimeter=0 $X=203925 $Y=116485 $dt=6
D21 11 5 p_dnw3 AREA=2.05478e-09 PJ=0 perimeter=0 $X=203925 $Y=135285 $dt=6
D22 11 5 p_dnw3 AREA=2.05478e-09 PJ=0 perimeter=0 $X=203925 $Y=154085 $dt=6
D23 11 5 p_dnw3 AREA=6.91743e-10 PJ=0 perimeter=0 $X=203925 $Y=172885 $dt=6
.ends dac6b_amp_n2
