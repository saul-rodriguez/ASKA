************************************************************************
* auCdl Netlist:
* 
* Library Name:  ASKA_REF_BIAS
* Top Cell Name: ref_bias
* View Name:     schematic
* Netlisted on:  Aug 26 08:30:29 2024
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.LDD
*.SCALE METER
.PARAM



************************************************************************
* Library Name: ASKA_REF_BIAS
* Cell Name:    ref_bias
* View Name:    schematic
************************************************************************

.SUBCKT ref_bias BIAS GNDA OUT1 OUT2 RES_BIAS VDDA VREF
*.PININFO BIAS:B GNDA:B OUT1:B OUT2:B RES_BIAS:B VDDA:B VREF:B
XM7 COM COM COM COM VDDA GNDA / ne3i_6 W=10u L=2u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ NRD=0.027 NRS=0.027 PD=2.096e-05 PS=2.096e-05 par1=4.0
XM12 net4 VREF COM COM VDDA GNDA / ne3i_6 W=10u L=2u M=14.0 AD=4.8e-12 
+ AS=4.8e-12 NRD=0.027 NRS=0.027 PD=2.096e-05 PS=2.096e-05 par1=14.0
XM24 net6 RES_BIAS COM COM VDDA GNDA / ne3i_6 W=10u L=2u M=14.0 AD=4.8e-12 
+ AS=4.8e-12 NRD=0.027 NRS=0.027 PD=2.096e-05 PS=2.096e-05 par1=14.0
MM10 GNDA GNDA GNDA GNDA NE3 W=10u L=5u M=5.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM9 BIAS BIAS net123 GNDA NE3 W=10u L=2u M=8.0 AD=2.7e-12 AS=3.225e-12 
+ PD=1.054e-05 PS=1.3145e-05 NRD=0.027 NRS=0.027
MM8 COM BIAS net5 GNDA NE3 W=10u L=2u M=8.0 AD=2.7e-12 AS=3.225e-12 
+ PD=1.054e-05 PS=1.3145e-05 NRD=0.027 NRS=0.027
MM26 net7 net123 GNDA GNDA NE3 W=10u L=5u M=1.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM13 net123 net123 GNDA GNDA NE3 W=10u L=5u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM25 net5 net123 GNDA GNDA NE3 W=10u L=5u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM6 VDDA VDDA VDDA VDDA PE3 W=10u L=2u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM5 VDDA VDDA VDDA VDDA PE3 W=10u L=10u M=4.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM28 net102 net102 VDDA VDDA PE3 W=10u L=2u M=2.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM0 net7 net7 net102 VDDA PE3 W=10u L=2u M=2.0 AD=2.7e-12 AS=4.8e-12 
+ PD=1.054e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM23 net6 net6 VDDA VDDA PE3 W=10u L=10u M=8.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM22 net4 net6 VDDA VDDA PE3 W=10u L=10u M=8.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM14 net8 net4 VDDA VDDA PE3 W=10u L=2u M=12.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM4 net1 net4 VDDA VDDA PE3 W=10u L=2u M=10.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM21 RES_BIAS net7 net8 VDDA PE3 W=10u L=1u M=12.0 AD=2.7e-12 AS=3.05e-12 
+ PD=1.054e-05 PS=1.22767e-05 NRD=0.027 NRS=0.027
MM3 OUT2 net7 net1 VDDA PE3 W=10u L=1u M=10.0 AD=2.7e-12 AS=3.12e-12 
+ PD=1.054e-05 PS=1.2624e-05 NRD=0.027 NRS=0.027
MM2 net2 net4 VDDA VDDA PE3 W=10u L=2u M=10.0 AD=4.8e-12 AS=4.8e-12 
+ PD=2.096e-05 PS=2.096e-05 NRD=0.027 NRS=0.027
MM1 OUT1 net7 net2 VDDA PE3 W=10u L=1u M=10.0 AD=2.7e-12 AS=3.12e-12 
+ PD=1.054e-05 PS=1.2624e-05 NRD=0.027 NRS=0.027
CC1 net4 net3 $[CMM5T] area=9e-10 perimeter=120.00000u M=8
RR0 net3 RES_BIAS 124.999K $SUB=GNDA $[RPP1K1_3] $W=4u $L=514.1u M=1
XC2 OUT2 GNDA GNDA / mosvc3 W=30u L=30u M=3.0 par1=3.0
XC0 OUT1 GNDA GNDA / mosvc3 W=30u L=30u M=3.0 par1=3.0
.ENDS


.SUBCKT mosvc3 G NW SB 
*.PININFO  G:B NW:B SB:B
.ENDS

.SUBCKT ne3i_6 D G S B NW SB 
*.PININFO  D:B G:B S:B B:B NW:B SB:B
.ENDS
