************************************************************************
* auCdl Netlist:
* 
* Library Name:  ALL_TESTS
* Top Cell Name: emir_test_1
* View Name:     schematic
* Netlisted on:  Jul 17 08:24:17 2024
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.LDD
*.SCALE METER
.PARAM



************************************************************************
* Library Name: ALL_TESTS
* Cell Name:    emir_test_1
* View Name:    schematic
************************************************************************

.SUBCKT emir_test_1 gnda vdda
*.PININFO gnda:B vdda:B
RR1 gnda vdda 1447.51 $[RPP1K1] $W=5u $L=25.0u M=1
RR0 gnda vdda 1447.51 $[RPP1K1] $W=5u $L=25.0u M=1
RR11 gnda vdda 1447.51 $[RPP1K1] $W=5u $L=25.0u M=1
.ENDS

