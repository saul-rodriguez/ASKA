* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : emir_test_2                                  *
* Netlisted  : Wed Aug  7 04:01:24 2024                     *
* PVS Version: 23.10-p043 Mon Oct 2 18:09:08 PDT 2023      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 R(rpp1k1) rpp1k1_2 p1trm(POS) p1trm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_CDNS_723017679630                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_CDNS_723017679630 2 3
** N=3 EP=2 FDC=1
R0 2 3 L=2.5e-05 W=5e-06 $[rpp1k1] $X=0 $Y=0 $dt=0
.ends rpp1k1_CDNS_723017679630

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: emir_test_2                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt emir_test_2 gnda vdda
** N=4 EP=2 FDC=7
X8 gnda vdda rpp1k1_CDNS_723017679630 $T=314165 13865 0 180 $X=288225 $Y=8645
X9 gnda vdda rpp1k1_CDNS_723017679630 $T=314165 23360 0 180 $X=288225 $Y=18140
X10 gnda vdda rpp1k1_CDNS_723017679630 $T=314165 34615 0 180 $X=288225 $Y=29395
X11 vdda gnda rpp1k1_CDNS_723017679630 $T=290815 57190 0 0 $X=289875 $Y=56970
X12 vdda gnda rpp1k1_CDNS_723017679630 $T=290815 65265 0 0 $X=289875 $Y=65045
X13 vdda gnda rpp1k1_CDNS_723017679630 $T=290815 72930 0 0 $X=289875 $Y=72710
X14 vdda gnda rpp1k1_CDNS_723017679630 $T=290815 80325 0 0 $X=289875 $Y=80105
.ends emir_test_2
