* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : bias                                         *
* Netlisted  : Mon Aug 26 08:37:01 2024                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(ne3) nem ndiff(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 1 MP(pe3) pem pdiff(D) p1trm(G) pdiff(S) nwtrm(B)
*.DEVTMPLT 2 NE3I_6() nemi_6 ndiff(D) p1trm(G) ndiff(S) pwitrm(B) dnwtrm(NW) bulk(SB)
*.DEVTMPLT 3 MOSVC3() mosvcm p1trm(G) nwtrm(NW) bulk(SB)
*.DEVTMPLT 4 Q(qpvc3) qpvmc bulk(C) nwtrm(B) pdiff(E)
*.DEVTMPLT 5 D(p_dnw) p_dnw bulk(POS) nwtrm(NEG)
*.DEVTMPLT 6 D(p_ddnw) p_ddnw bulk(POS) dnwtrm(NEG)
*.DEVTMPLT 7 D(p_dipdnwmv) p_dipwmv pwitrm(POS) dnwtrm(NEG)
*.DEVTMPLT 8 D(p_dnw3) p_dnwm bulk(POS) nwtrm(NEG)
*.DEVTMPLT 9 R(rpp1k1_3) rpp1k1_s p1trm(POS) p1trm(NEG) bulk(SUB)
*.DEVTMPLT 10 R(rpp1k1_3) rpp1k1_n p1trm(POS) p1trm(NEG) nwtrm(SUB)
*.DEVTMPLT 11 C(cmm5t) cmim capm(POS) m4trm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NE3I_6                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NE3I_6 D G S B NW SB
.ends NE3I_6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MOSVC3                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MOSVC3 G NW SB
.ends MOSVC3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724654214590                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724654214590 1 2 3 4 5
** N=5 EP=5 FDC=11
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=1
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=1
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=1
M4 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=6160 $Y=0 $dt=1
M5 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7700 $Y=0 $dt=1
M6 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=9240 $Y=0 $dt=1
M7 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10780 $Y=0 $dt=1
M8 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12320 $Y=0 $dt=1
M9 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=13860 $Y=0 $dt=1
D10 5 4 p_dnw3 AREA=2.15633e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=8
.ends pe3_CDNS_724654214590

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724654214591                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724654214591 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 ne3 L=5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
.ends ne3_CDNS_724654214591

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724654214592                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724654214592 1 2 3 4 5
** N=5 EP=5 FDC=13
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=1
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=1
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=1
M4 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=6160 $Y=0 $dt=1
M5 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7700 $Y=0 $dt=1
M6 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=9240 $Y=0 $dt=1
M7 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10780 $Y=0 $dt=1
M8 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12320 $Y=0 $dt=1
M9 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=13860 $Y=0 $dt=1
M10 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=15400 $Y=0 $dt=1
M11 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=16940 $Y=0 $dt=1
D12 5 4 p_dnw3 AREA=2.52778e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=8
.ends pe3_CDNS_724654214592

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724654214593                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724654214593 1 2 3 4
** N=4 EP=4 FDC=3
M0 2 2 1 3 pe3 L=2e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 2 3 pe3 L=2e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=2540 $Y=0 $dt=1
D2 4 3 p_dnw3 AREA=9.11736e-11 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=8
.ends pe3_CDNS_724654214593

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_724654214594                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_724654214594 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.0005141 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=9
.ends rpp1k1_3_CDNS_724654214594

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724654214595                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724654214595 1 2 3 4
** N=4 EP=4 FDC=8
M0 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
M1 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=2540 $Y=0 $dt=0
M2 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=5080 $Y=0 $dt=0
M3 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=7620 $Y=0 $dt=0
M4 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=10160 $Y=0 $dt=0
M5 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=12700 $Y=0 $dt=0
M6 3 2 1 4 ne3 L=2e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=15240 $Y=0 $dt=0
M7 1 2 3 4 ne3 L=2e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=17780 $Y=0 $dt=0
.ends ne3_CDNS_724654214595

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724654214599                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724654214599 1 2 3
*.DEVICECLIMB
** N=4 EP=3 FDC=1
M0 3 2 1 1 pe3 L=2e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_724654214599

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246542145910                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246542145910 1 2 3
*.DEVICECLIMB
** N=4 EP=3 FDC=1
M0 3 2 1 1 pe3 L=1e-05 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_7246542145910

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3i_6_CDNS_724654214598                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3i_6_CDNS_724654214598 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=1
X0 1 2 3 1 4 5 NE3I_6 w=1e-05 l=2e-06 as=4.8e-12 ad=4.8e-12 ps=2.096e-05 pd=2.096e-05 $X=0 $Y=0 $dt=2
.ends ne3i_6_CDNS_724654214598

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A3                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A3 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=2
X0 1 4 5 6 7 ne3i_6_CDNS_724654214598 $T=4060 14570 1 0 $X=0 $Y=0
X1 1 2 3 6 7 ne3i_6_CDNS_724654214598 $T=7460 14570 1 0 $X=3400 $Y=0
.ends MASCO__A3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A4                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A4 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=2
X0 1 4 5 6 7 ne3i_6_CDNS_724654214598 $T=4060 4450 0 0 $X=0 $Y=0
X1 1 2 3 6 7 ne3i_6_CDNS_724654214598 $T=7460 4450 0 0 $X=3400 $Y=0
.ends MASCO__A4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__B5                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__B5 1 2 3 4 5 6 7 8 9 10
+ 11
*.DEVICECLIMB
** N=11 EP=11 FDC=4
X0 1 10 6 5 3 2 11 MASCO__A3 $T=0 14680 0 0 $X=0 $Y=14680
X1 1 8 7 9 4 2 11 MASCO__A4 $T=0 0 0 0 $X=0 $Y=0
.ends MASCO__B5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ref_bias                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ref_bias GNDA VDDA BIAS RES_BIAS OUT2 OUT1 VREF
** N=18 EP=7 FDC=187
X556 14 8 OUT1 VDDA GNDA pe3_CDNS_724654214590 $T=189280 150320 0 0 $X=187770 $Y=149290
X557 15 8 OUT2 VDDA GNDA pe3_CDNS_724654214590 $T=213190 150320 0 0 $X=211680 $Y=149290
X558 GNDA GNDA GNDA ne3_CDNS_724654214591 $T=17980 14080 0 0 $X=17180 $Y=13680
X559 GNDA GNDA GNDA ne3_CDNS_724654214591 $T=17980 30170 0 0 $X=17180 $Y=29770
X560 GNDA 9 10 ne3_CDNS_724654214591 $T=24220 14080 0 0 $X=23420 $Y=13680
X561 GNDA 9 9 ne3_CDNS_724654214591 $T=24220 30170 0 0 $X=23420 $Y=29770
X562 GNDA 9 9 ne3_CDNS_724654214591 $T=30460 14080 0 0 $X=29660 $Y=13680
X563 GNDA 9 10 ne3_CDNS_724654214591 $T=30460 30170 0 0 $X=29660 $Y=29770
X564 GNDA 9 8 ne3_CDNS_724654214591 $T=36700 14080 0 0 $X=35900 $Y=13680
X565 GNDA 9 9 ne3_CDNS_724654214591 $T=36700 30170 0 0 $X=35900 $Y=29770
X566 GNDA 9 9 ne3_CDNS_724654214591 $T=42940 14080 0 0 $X=42140 $Y=13680
X567 GNDA 9 10 ne3_CDNS_724654214591 $T=42940 30170 0 0 $X=42140 $Y=29770
X568 GNDA 9 10 ne3_CDNS_724654214591 $T=49180 14080 0 0 $X=48380 $Y=13680
X569 GNDA GNDA GNDA ne3_CDNS_724654214591 $T=49180 30170 0 0 $X=48380 $Y=29770
X570 GNDA GNDA GNDA ne3_CDNS_724654214591 $T=55420 14080 0 0 $X=54620 $Y=13680
X571 GNDA GNDA GNDA ne3_CDNS_724654214591 $T=55420 30170 0 0 $X=54620 $Y=29770
X572 13 8 RES_BIAS VDDA GNDA pe3_CDNS_724654214592 $T=162340 150320 0 0 $X=160830 $Y=149290
X573 VDDA 12 VDDA GNDA pe3_CDNS_724654214593 $T=138060 190125 0 0 $X=136550 $Y=189095
X574 12 8 VDDA GNDA pe3_CDNS_724654214593 $T=147620 190125 0 0 $X=146110 $Y=189095
X575 RES_BIAS 18 GNDA rpp1k1_3_CDNS_724654214594 $T=87870 117335 0 0 $X=82710 $Y=117115
X576 9 BIAS BIAS GNDA ne3_CDNS_724654214595 $T=17545 54415 0 0 $X=16745 $Y=54015
X577 10 BIAS 11 GNDA ne3_CDNS_724654214595 $T=42480 54195 0 0 $X=41680 $Y=53795
X578 VDDA VDDA VDDA pe3_CDNS_724654214599 $T=165675 175935 0 0 $X=164165 $Y=174905
X579 VDDA VDDA VDDA pe3_CDNS_724654214599 $T=165675 195955 0 0 $X=164165 $Y=194925
X580 VDDA 17 14 pe3_CDNS_724654214599 $T=168915 175935 0 0 $X=167405 $Y=174905
X581 VDDA 17 15 pe3_CDNS_724654214599 $T=168915 195955 0 0 $X=167405 $Y=194925
X582 VDDA 17 15 pe3_CDNS_724654214599 $T=172155 175935 0 0 $X=170645 $Y=174905
X583 VDDA 17 13 pe3_CDNS_724654214599 $T=172155 195955 0 0 $X=170645 $Y=194925
X584 VDDA 17 13 pe3_CDNS_724654214599 $T=175395 175935 0 0 $X=173885 $Y=174905
X585 VDDA 17 14 pe3_CDNS_724654214599 $T=175395 195955 0 0 $X=173885 $Y=194925
X586 VDDA 17 14 pe3_CDNS_724654214599 $T=178635 175935 0 0 $X=177125 $Y=174905
X587 VDDA 17 15 pe3_CDNS_724654214599 $T=178635 195955 0 0 $X=177125 $Y=194925
X588 VDDA 17 13 pe3_CDNS_724654214599 $T=181875 175935 0 0 $X=180365 $Y=174905
X589 VDDA 17 15 pe3_CDNS_724654214599 $T=181875 195955 0 0 $X=180365 $Y=194925
X590 VDDA 17 15 pe3_CDNS_724654214599 $T=185115 175935 0 0 $X=183605 $Y=174905
X591 VDDA 17 13 pe3_CDNS_724654214599 $T=185115 195955 0 0 $X=183605 $Y=194925
X592 VDDA 17 13 pe3_CDNS_724654214599 $T=188355 175935 0 0 $X=186845 $Y=174905
X593 VDDA 17 14 pe3_CDNS_724654214599 $T=188355 195955 0 0 $X=186845 $Y=194925
X594 VDDA 17 14 pe3_CDNS_724654214599 $T=191595 175935 0 0 $X=190085 $Y=174905
X595 VDDA 17 13 pe3_CDNS_724654214599 $T=191595 195955 0 0 $X=190085 $Y=194925
X596 VDDA 17 13 pe3_CDNS_724654214599 $T=194835 175935 0 0 $X=193325 $Y=174905
X597 VDDA 17 15 pe3_CDNS_724654214599 $T=194835 195955 0 0 $X=193325 $Y=194925
X598 VDDA 17 15 pe3_CDNS_724654214599 $T=198075 175935 0 0 $X=196565 $Y=174905
X599 VDDA 17 13 pe3_CDNS_724654214599 $T=198075 195955 0 0 $X=196565 $Y=194925
X600 VDDA 17 13 pe3_CDNS_724654214599 $T=201315 175935 0 0 $X=199805 $Y=174905
X601 VDDA 17 14 pe3_CDNS_724654214599 $T=201315 195955 0 0 $X=199805 $Y=194925
X602 VDDA 17 14 pe3_CDNS_724654214599 $T=204555 175935 0 0 $X=203045 $Y=174905
X603 VDDA 17 13 pe3_CDNS_724654214599 $T=204555 195955 0 0 $X=203045 $Y=194925
X604 VDDA 17 14 pe3_CDNS_724654214599 $T=207795 175935 0 0 $X=206285 $Y=174905
X605 VDDA 17 15 pe3_CDNS_724654214599 $T=207795 195955 0 0 $X=206285 $Y=194925
X606 VDDA 17 15 pe3_CDNS_724654214599 $T=211035 175935 0 0 $X=209525 $Y=174905
X607 VDDA 17 13 pe3_CDNS_724654214599 $T=211035 195955 0 0 $X=209525 $Y=194925
X608 VDDA 17 13 pe3_CDNS_724654214599 $T=214275 175935 0 0 $X=212765 $Y=174905
X609 VDDA 17 14 pe3_CDNS_724654214599 $T=214275 195955 0 0 $X=212765 $Y=194925
X610 VDDA 17 14 pe3_CDNS_724654214599 $T=217515 175935 0 0 $X=216005 $Y=174905
X611 VDDA 17 15 pe3_CDNS_724654214599 $T=217515 195955 0 0 $X=216005 $Y=194925
X612 VDDA VDDA VDDA pe3_CDNS_724654214599 $T=220755 175935 0 0 $X=219245 $Y=174905
X613 VDDA VDDA VDDA pe3_CDNS_724654214599 $T=220755 195955 0 0 $X=219245 $Y=194925
X614 VDDA VDDA VDDA pe3_CDNS_7246542145910 $T=12010 172320 0 0 $X=10500 $Y=171290
X615 VDDA VDDA VDDA pe3_CDNS_7246542145910 $T=12010 190000 0 0 $X=10500 $Y=188970
X616 VDDA 16 16 pe3_CDNS_7246542145910 $T=23250 172320 0 0 $X=21740 $Y=171290
X617 VDDA 16 17 pe3_CDNS_7246542145910 $T=23250 190000 0 0 $X=21740 $Y=188970
X618 VDDA 16 17 pe3_CDNS_7246542145910 $T=34490 172320 0 0 $X=32980 $Y=171290
X619 VDDA 16 16 pe3_CDNS_7246542145910 $T=34490 190000 0 0 $X=32980 $Y=188970
X620 VDDA 16 16 pe3_CDNS_7246542145910 $T=45730 172320 0 0 $X=44220 $Y=171290
X621 VDDA 16 17 pe3_CDNS_7246542145910 $T=45730 190000 0 0 $X=44220 $Y=188970
X622 VDDA 16 17 pe3_CDNS_7246542145910 $T=56970 172320 0 0 $X=55460 $Y=171290
X623 VDDA 16 16 pe3_CDNS_7246542145910 $T=56970 190000 0 0 $X=55460 $Y=188970
X624 VDDA 16 16 pe3_CDNS_7246542145910 $T=68210 172320 0 0 $X=66700 $Y=171290
X625 VDDA 16 17 pe3_CDNS_7246542145910 $T=68210 190000 0 0 $X=66700 $Y=188970
X626 VDDA 16 17 pe3_CDNS_7246542145910 $T=79450 172320 0 0 $X=77940 $Y=171290
X627 VDDA 16 16 pe3_CDNS_7246542145910 $T=79450 190000 0 0 $X=77940 $Y=188970
X628 VDDA 16 16 pe3_CDNS_7246542145910 $T=90690 172320 0 0 $X=89180 $Y=171290
X629 VDDA 16 17 pe3_CDNS_7246542145910 $T=90690 190000 0 0 $X=89180 $Y=188970
X630 VDDA 16 17 pe3_CDNS_7246542145910 $T=101930 172320 0 0 $X=100420 $Y=171290
X631 VDDA 16 16 pe3_CDNS_7246542145910 $T=101930 190000 0 0 $X=100420 $Y=188970
X632 VDDA VDDA VDDA pe3_CDNS_7246542145910 $T=113170 172320 0 0 $X=111660 $Y=171290
X633 VDDA VDDA VDDA pe3_CDNS_7246542145910 $T=113170 190000 0 0 $X=111660 $Y=188970
X634 11 VDDA 11 11 11 17 16 RES_BIAS 11 VREF
+ GNDA MASCO__B5 $T=9330 114030 0 0 $X=9330 $Y=114030
X635 11 VDDA 16 17 RES_BIAS 17 16 RES_BIAS VREF VREF
+ GNDA MASCO__B5 $T=16130 114030 0 0 $X=16130 $Y=114030
X636 11 VDDA 16 17 RES_BIAS 17 16 RES_BIAS VREF VREF
+ GNDA MASCO__B5 $T=22930 114030 0 0 $X=22930 $Y=114030
X637 11 VDDA 16 17 RES_BIAS 17 16 RES_BIAS VREF VREF
+ GNDA MASCO__B5 $T=29730 114030 0 0 $X=29730 $Y=114030
X638 11 VDDA 16 17 RES_BIAS 17 16 RES_BIAS VREF VREF
+ GNDA MASCO__B5 $T=36530 114030 0 0 $X=36530 $Y=114030
X639 11 VDDA 16 17 RES_BIAS 17 16 RES_BIAS VREF VREF
+ GNDA MASCO__B5 $T=43330 114030 0 0 $X=43330 $Y=114030
X640 11 VDDA 16 17 RES_BIAS 17 16 RES_BIAS VREF VREF
+ GNDA MASCO__B5 $T=50130 114030 0 0 $X=50130 $Y=114030
X641 11 VDDA 16 17 RES_BIAS 11 11 11 VREF 11
+ GNDA MASCO__B5 $T=56930 114030 0 0 $X=56930 $Y=114030
X642 OUT2 GNDA GNDA MOSVC3 w=3e-05 l=3e-05 $X=85530 $Y=8110 $dt=3
X643 OUT2 GNDA GNDA MOSVC3 w=3e-05 l=3e-05 $X=85530 $Y=39350 $dt=3
X644 OUT2 GNDA GNDA MOSVC3 w=3e-05 l=3e-05 $X=85530 $Y=70590 $dt=3
X645 OUT1 GNDA GNDA MOSVC3 w=3e-05 l=3e-05 $X=122495 $Y=8050 $dt=3
X646 OUT1 GNDA GNDA MOSVC3 w=3e-05 l=3e-05 $X=122495 $Y=39290 $dt=3
X647 OUT1 GNDA GNDA MOSVC3 w=3e-05 l=3e-05 $X=122495 $Y=70530 $dt=3
D6 GNDA VDDA p_dnw AREA=2.36318e-09 PJ=0.00033402 perimeter=0.00033402 $X=4385 $Y=163650 $dt=5
D7 GNDA VDDA p_dnw AREA=2.57209e-10 PJ=8.388e-05 perimeter=8.388e-05 $X=134410 $Y=183535 $dt=5
D8 GNDA VDDA p_dnw AREA=1.81014e-09 PJ=0.00023539 perimeter=0.00023539 $X=158410 $Y=166295 $dt=5
D9 GNDA VDDA p_dnw AREA=8.15582e-10 PJ=0.0001871 perimeter=0.0001871 $X=158690 $Y=143730 $dt=5
D10 GNDA VDDA p_dnw AREA=9.45702e-09 PJ=0.00040696 perimeter=0.00040696 $X=159475 $Y=6005 $dt=5
D11 GNDA VDDA p_ddnw AREA=1.66704e-09 PJ=0.0001998 perimeter=0.0001998 $X=8060 $Y=112760 $dt=6
D12 11 VDDA p_dipdnwmv AREA=9.57098e-10 PJ=0.000169 perimeter=0.000169 $X=11910 $Y=116610 $dt=7
D13 GNDA VDDA p_dnw3 AREA=1.37701e-09 PJ=0 perimeter=0 $X=10500 $Y=171290 $dt=8
D14 GNDA VDDA p_dnw3 AREA=1.37701e-09 PJ=0 perimeter=0 $X=10500 $Y=188970 $dt=8
D15 GNDA GNDA p_dnw3 AREA=2.03309e-10 PJ=0.00024988 perimeter=0.00024988 $X=85100 $Y=7310 $dt=8
D16 GNDA GNDA p_dnw3 AREA=2.03309e-10 PJ=0.00024988 perimeter=0.00024988 $X=122065 $Y=7250 $dt=8
D17 GNDA VDDA p_dnw3 AREA=7.24806e-10 PJ=0 perimeter=0 $X=164165 $Y=174905 $dt=8
D18 GNDA VDDA p_dnw3 AREA=7.24806e-10 PJ=0 perimeter=0 $X=164165 $Y=194925 $dt=8
C19 17 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=161615 $Y=8145 $dt=11
C20 17 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=161615 $Y=39745 $dt=11
C21 17 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=161615 $Y=71345 $dt=11
C22 17 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=161615 $Y=102945 $dt=11
C23 17 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=196615 $Y=8145 $dt=11
C24 17 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=196615 $Y=39745 $dt=11
C25 17 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=196615 $Y=71345 $dt=11
C26 17 18 area=9e-10 perimeter=0.00012 $[cmm5t] $X=196615 $Y=102945 $dt=11
.ends ref_bias

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246542145911                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246542145911 1 2 3 4 5
** N=5 EP=5 FDC=5
M0 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=1
M2 3 2 1 4 pe3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=1
M3 1 2 3 4 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=1
D4 5 4 p_dnw3 AREA=1.04198e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=8
.ends pe3_CDNS_7246542145911

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7246542145912                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7246542145912 1 2 3 4
** N=4 EP=4 FDC=4
M0 3 2 1 4 ne3 L=1e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
M1 1 2 3 4 ne3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=1540 $Y=0 $dt=0
M2 3 2 1 4 ne3 L=1e-06 W=1e-05 AD=2.7e-12 AS=2.7e-12 PD=1.054e-05 PS=1.054e-05 $X=3080 $Y=0 $dt=0
M3 1 2 3 4 ne3 L=1e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=4620 $Y=0 $dt=0
.ends ne3_CDNS_7246542145912

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7246542145913                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7246542145913 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.0005215 W=8e-06 $[rpp1k1_3] $SUB=3 $X=-8220 $Y=0 $dt=9
.ends rpp1k1_3_CDNS_7246542145913

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7246542145914                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7246542145914 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.00082283 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=9
.ends rpp1k1_3_CDNS_7246542145914

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7246542145915                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7246542145915 1 2 3 4
** N=4 EP=4 FDC=1
M0 3 2 1 4 ne3 L=1e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
.ends ne3_CDNS_7246542145915

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246542145916                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246542145916 1 2 3 4
*.DEVICECLIMB
** N=5 EP=4 FDC=1
M0 3 2 1 4 pe3 L=5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_7246542145916

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246542145917                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246542145917 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 3 2 1 4 pe3 L=5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
D1 5 4 p_dnw3 AREA=9.67212e-11 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=8
.ends pe3_CDNS_7246542145917

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7246542145918                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7246542145918 1 2 3
** N=3 EP=3 FDC=1
M0 2 2 1 3 ne3 L=2e-06 W=1e-06 AD=4.8e-13 AS=4.8e-13 PD=2.96e-06 PS=2.96e-06 $X=0 $Y=0 $dt=0
.ends ne3_CDNS_7246542145918

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246542145919                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246542145919 1 2 3
*.DEVICECLIMB
** N=4 EP=3 FDC=1
M0 3 2 1 1 pe3 L=1e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_7246542145919

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7246542145920                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7246542145920 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.00082283 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=9
.ends rpp1k1_3_CDNS_7246542145920

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: bandgap_su                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt bandgap_su GNDA VDD3A BIAS OUT
** N=24 EP=4 FDC=165
X308 GNDA GNDA GNDA ne3_CDNS_724654214591 $T=44780 15300 0 0 $X=43980 $Y=14900
X309 GNDA GNDA GNDA ne3_CDNS_724654214591 $T=44780 37440 1 0 $X=43980 $Y=26870
X310 GNDA 11 11 ne3_CDNS_724654214591 $T=51020 15300 0 0 $X=50220 $Y=14900
X311 GNDA 11 14 ne3_CDNS_724654214591 $T=51020 37440 1 0 $X=50220 $Y=26870
X312 GNDA 11 14 ne3_CDNS_724654214591 $T=57260 15300 0 0 $X=56460 $Y=14900
X313 GNDA 11 11 ne3_CDNS_724654214591 $T=57260 37440 1 0 $X=56460 $Y=26870
X314 GNDA 11 11 ne3_CDNS_724654214591 $T=63500 15300 0 0 $X=62700 $Y=14900
X315 GNDA 11 14 ne3_CDNS_724654214591 $T=63500 37440 1 0 $X=62700 $Y=26870
X316 GNDA 11 14 ne3_CDNS_724654214591 $T=69740 15300 0 0 $X=68940 $Y=14900
X317 GNDA 11 11 ne3_CDNS_724654214591 $T=69740 37440 1 0 $X=68940 $Y=26870
X318 GNDA 11 11 ne3_CDNS_724654214591 $T=75980 15300 0 0 $X=75180 $Y=14900
X319 GNDA 11 14 ne3_CDNS_724654214591 $T=75980 37440 1 0 $X=75180 $Y=26870
X320 GNDA 11 14 ne3_CDNS_724654214591 $T=82220 15300 0 0 $X=81420 $Y=14900
X321 GNDA 11 11 ne3_CDNS_724654214591 $T=82220 37440 1 0 $X=81420 $Y=26870
X322 GNDA 11 11 ne3_CDNS_724654214591 $T=88460 15300 0 0 $X=87660 $Y=14900
X323 GNDA 11 14 ne3_CDNS_724654214591 $T=88460 37440 1 0 $X=87660 $Y=26870
X324 GNDA 11 14 ne3_CDNS_724654214591 $T=94700 15300 0 0 $X=93900 $Y=14900
X325 GNDA 11 11 ne3_CDNS_724654214591 $T=94700 37440 1 0 $X=93900 $Y=26870
X326 GNDA GNDA GNDA ne3_CDNS_724654214591 $T=100940 15300 0 0 $X=100140 $Y=14900
X327 GNDA GNDA GNDA ne3_CDNS_724654214591 $T=100940 37440 1 0 $X=100140 $Y=26870
X380 8 6 6 VDD3A GNDA pe3_CDNS_7246542145911 $T=9635 78185 0 0 $X=8125 $Y=77155
X381 5 6 19 VDD3A GNDA pe3_CDNS_7246542145911 $T=23440 78185 0 0 $X=21930 $Y=77155
X382 7 BIAS BIAS GNDA ne3_CDNS_7246542145912 $T=10345 55405 0 0 $X=9545 $Y=55005
X383 16 BIAS 6 GNDA ne3_CDNS_7246542145912 $T=22730 55545 0 0 $X=21930 $Y=55145
X384 GNDA 14 OUT GNDA ne3_CDNS_7246542145912 $T=95790 103175 0 0 $X=94990 $Y=102775
X385 9 21 GNDA rpp1k1_3_CDNS_7246542145913 $T=287735 7255 1 180 $X=159445 $Y=7035
X386 OUT 22 GNDA rpp1k1_3_CDNS_7246542145914 $T=123895 47740 0 0 $X=118735 $Y=47520
X387 GNDA GNDA GNDA GNDA ne3_CDNS_7246542145915 $T=13130 16755 0 0 $X=12330 $Y=16355
X388 GNDA GNDA GNDA GNDA ne3_CDNS_7246542145915 $T=13130 38815 1 0 $X=12330 $Y=28245
X389 GNDA 7 16 GNDA ne3_CDNS_7246542145915 $T=15370 16755 0 0 $X=14570 $Y=16355
X390 GNDA 7 7 GNDA ne3_CDNS_7246542145915 $T=15370 38815 1 0 $X=14570 $Y=28245
X391 GNDA 7 7 GNDA ne3_CDNS_7246542145915 $T=17610 16755 0 0 $X=16810 $Y=16355
X392 GNDA 7 16 GNDA ne3_CDNS_7246542145915 $T=17610 38815 1 0 $X=16810 $Y=28245
X393 GNDA 7 17 GNDA ne3_CDNS_7246542145915 $T=19850 16755 0 0 $X=19050 $Y=16355
X394 GNDA 7 18 GNDA ne3_CDNS_7246542145915 $T=19850 38815 1 0 $X=19050 $Y=28245
X395 GNDA 7 16 GNDA ne3_CDNS_7246542145915 $T=22090 16755 0 0 $X=21290 $Y=16355
X396 GNDA 7 7 GNDA ne3_CDNS_7246542145915 $T=22090 38815 1 0 $X=21290 $Y=28245
X397 GNDA 7 7 GNDA ne3_CDNS_7246542145915 $T=24330 16755 0 0 $X=23530 $Y=16355
X398 GNDA 7 16 GNDA ne3_CDNS_7246542145915 $T=24330 38815 1 0 $X=23530 $Y=28245
X399 GNDA GNDA GNDA GNDA ne3_CDNS_7246542145915 $T=26570 16755 0 0 $X=25770 $Y=16355
X400 GNDA GNDA GNDA GNDA ne3_CDNS_7246542145915 $T=26570 38815 1 0 $X=25770 $Y=28245
X401 17 OUT 13 GNDA ne3_CDNS_7246542145915 $T=97960 125180 0 0 $X=97160 $Y=124780
X402 17 15 20 GNDA ne3_CDNS_7246542145915 $T=100200 125180 0 0 $X=99400 $Y=124780
X403 19 19 19 VDD3A pe3_CDNS_7246542145916 $T=43105 60145 0 0 $X=41595 $Y=59115
X404 19 19 19 VDD3A pe3_CDNS_7246542145916 $T=43105 83765 1 0 $X=41595 $Y=72735
X405 19 10 14 VDD3A pe3_CDNS_7246542145916 $T=49345 60145 0 0 $X=47835 $Y=59115
X406 19 9 11 VDD3A pe3_CDNS_7246542145916 $T=49345 83765 1 0 $X=47835 $Y=72735
X407 19 9 11 VDD3A pe3_CDNS_7246542145916 $T=55585 60145 0 0 $X=54075 $Y=59115
X408 19 10 14 VDD3A pe3_CDNS_7246542145916 $T=55585 83765 1 0 $X=54075 $Y=72735
X409 VDD3A 12 12 VDD3A pe3_CDNS_7246542145916 $T=59655 129400 1 0 $X=58145 $Y=118370
X410 19 10 14 VDD3A pe3_CDNS_7246542145916 $T=61825 60145 0 0 $X=60315 $Y=59115
X411 19 9 11 VDD3A pe3_CDNS_7246542145916 $T=61825 83765 1 0 $X=60315 $Y=72735
X412 VDD3A 12 10 VDD3A pe3_CDNS_7246542145916 $T=65895 129400 1 0 $X=64385 $Y=118370
X413 19 9 11 VDD3A pe3_CDNS_7246542145916 $T=68065 60145 0 0 $X=66555 $Y=59115
X414 19 10 14 VDD3A pe3_CDNS_7246542145916 $T=68065 83765 1 0 $X=66555 $Y=72735
X415 19 10 14 VDD3A pe3_CDNS_7246542145916 $T=74305 60145 0 0 $X=72795 $Y=59115
X416 19 9 11 VDD3A pe3_CDNS_7246542145916 $T=74305 83765 1 0 $X=72795 $Y=72735
X417 VDD3A 13 13 VDD3A pe3_CDNS_7246542145916 $T=79075 125320 0 0 $X=77565 $Y=124290
X418 19 9 11 VDD3A pe3_CDNS_7246542145916 $T=80545 60145 0 0 $X=79035 $Y=59115
X419 19 10 14 VDD3A pe3_CDNS_7246542145916 $T=80545 83765 1 0 $X=79035 $Y=72735
X420 VDD3A 13 20 VDD3A pe3_CDNS_7246542145916 $T=85315 125320 0 0 $X=83805 $Y=124290
X421 19 10 14 VDD3A pe3_CDNS_7246542145916 $T=86785 60145 0 0 $X=85275 $Y=59115
X422 19 9 11 VDD3A pe3_CDNS_7246542145916 $T=86785 83765 1 0 $X=85275 $Y=72735
X423 19 9 11 VDD3A pe3_CDNS_7246542145916 $T=93025 60145 0 0 $X=91515 $Y=59115
X424 19 10 14 VDD3A pe3_CDNS_7246542145916 $T=93025 83765 1 0 $X=91515 $Y=72735
X425 19 19 19 VDD3A pe3_CDNS_7246542145916 $T=99265 60145 0 0 $X=97755 $Y=59115
X426 19 19 19 VDD3A pe3_CDNS_7246542145916 $T=99265 83765 1 0 $X=97755 $Y=72735
X427 12 20 18 VDD3A GNDA pe3_CDNS_7246542145917 $T=62750 104210 0 0 $X=61240 $Y=103180
X428 GNDA 15 GNDA ne3_CDNS_7246542145918 $T=110195 126990 0 0 $X=109395 $Y=126590
X429 15 23 GNDA ne3_CDNS_7246542145918 $T=110195 130510 0 0 $X=109395 $Y=130110
X430 23 VDD3A GNDA ne3_CDNS_7246542145918 $T=110195 134045 0 0 $X=109395 $Y=133645
X431 VDD3A VDD3A VDD3A pe3_CDNS_7246542145919 $T=10660 106140 0 0 $X=9150 $Y=105110
X432 VDD3A VDD3A VDD3A pe3_CDNS_7246542145919 $T=10660 129120 1 0 $X=9150 $Y=118090
X433 VDD3A 8 OUT pe3_CDNS_7246542145919 $T=12900 106140 0 0 $X=11390 $Y=105110
X434 VDD3A 8 OUT pe3_CDNS_7246542145919 $T=12900 129120 1 0 $X=11390 $Y=118090
X435 VDD3A 8 OUT pe3_CDNS_7246542145919 $T=15140 106140 0 0 $X=13630 $Y=105110
X436 VDD3A 8 OUT pe3_CDNS_7246542145919 $T=15140 129120 1 0 $X=13630 $Y=118090
X437 VDD3A 8 5 pe3_CDNS_7246542145919 $T=17380 106140 0 0 $X=15870 $Y=105110
X438 VDD3A 8 8 pe3_CDNS_7246542145919 $T=17380 129120 1 0 $X=15870 $Y=118090
X439 VDD3A 8 OUT pe3_CDNS_7246542145919 $T=19620 106140 0 0 $X=18110 $Y=105110
X440 VDD3A 8 OUT pe3_CDNS_7246542145919 $T=19620 129120 1 0 $X=18110 $Y=118090
X441 VDD3A 8 OUT pe3_CDNS_7246542145919 $T=21860 106140 0 0 $X=20350 $Y=105110
X442 VDD3A 8 OUT pe3_CDNS_7246542145919 $T=21860 129120 1 0 $X=20350 $Y=118090
X443 VDD3A 8 8 pe3_CDNS_7246542145919 $T=24100 106140 0 0 $X=22590 $Y=105110
X444 VDD3A 8 5 pe3_CDNS_7246542145919 $T=24100 129120 1 0 $X=22590 $Y=118090
X445 VDD3A 8 5 pe3_CDNS_7246542145919 $T=26340 106140 0 0 $X=24830 $Y=105110
X446 VDD3A 8 8 pe3_CDNS_7246542145919 $T=26340 129120 1 0 $X=24830 $Y=118090
X447 VDD3A 8 OUT pe3_CDNS_7246542145919 $T=28580 106140 0 0 $X=27070 $Y=105110
X448 VDD3A 8 OUT pe3_CDNS_7246542145919 $T=28580 129120 1 0 $X=27070 $Y=118090
X449 VDD3A 8 OUT pe3_CDNS_7246542145919 $T=30820 106140 0 0 $X=29310 $Y=105110
X450 VDD3A 8 OUT pe3_CDNS_7246542145919 $T=30820 129120 1 0 $X=29310 $Y=118090
X451 VDD3A 8 8 pe3_CDNS_7246542145919 $T=33060 106140 0 0 $X=31550 $Y=105110
X452 VDD3A 8 5 pe3_CDNS_7246542145919 $T=33060 129120 1 0 $X=31550 $Y=118090
X453 VDD3A 8 OUT pe3_CDNS_7246542145919 $T=35300 106140 0 0 $X=33790 $Y=105110
X454 VDD3A 8 OUT pe3_CDNS_7246542145919 $T=35300 129120 1 0 $X=33790 $Y=118090
X455 VDD3A 8 OUT pe3_CDNS_7246542145919 $T=37540 106140 0 0 $X=36030 $Y=105110
X456 VDD3A 8 OUT pe3_CDNS_7246542145919 $T=37540 129120 1 0 $X=36030 $Y=118090
X457 VDD3A VDD3A VDD3A pe3_CDNS_7246542145919 $T=39780 106140 0 0 $X=38270 $Y=105110
X458 VDD3A VDD3A VDD3A pe3_CDNS_7246542145919 $T=39780 129120 1 0 $X=38270 $Y=118090
X459 OUT 24 GNDA rpp1k1_3_CDNS_7246542145920 $T=123895 96235 0 0 $X=118735 $Y=96015
X460 22 9 GNDA rpp1k1_3_CDNS_7246542145920 $T=213685 47740 0 0 $X=208525 $Y=47520
X461 24 10 GNDA rpp1k1_3_CDNS_7246542145920 $T=213685 96235 0 0 $X=208525 $Y=96015
Q0 GNDA GNDA 21 qpvc3 $X=302595 $Y=9520 $dt=4
Q1 GNDA GNDA 21 qpvc3 $X=302595 $Y=26270 $dt=4
Q2 GNDA GNDA 21 qpvc3 $X=302595 $Y=43020 $dt=4
Q3 GNDA GNDA 21 qpvc3 $X=302595 $Y=59770 $dt=4
Q4 GNDA GNDA 21 qpvc3 $X=302595 $Y=76520 $dt=4
Q5 GNDA GNDA 21 qpvc3 $X=302595 $Y=93270 $dt=4
Q6 GNDA GNDA 21 qpvc3 $X=302595 $Y=110020 $dt=4
Q7 GNDA GNDA 21 qpvc3 $X=302595 $Y=126770 $dt=4
Q8 GNDA GNDA 21 qpvc3 $X=319350 $Y=9520 $dt=4
Q9 GNDA GNDA 21 qpvc3 $X=319350 $Y=26270 $dt=4
Q10 GNDA GNDA 21 qpvc3 $X=319350 $Y=43020 $dt=4
Q11 GNDA GNDA 10 qpvc3 $X=319350 $Y=59770 $dt=4
Q12 GNDA GNDA 21 qpvc3 $X=319350 $Y=76520 $dt=4
Q13 GNDA GNDA 21 qpvc3 $X=319350 $Y=93270 $dt=4
Q14 GNDA GNDA 21 qpvc3 $X=319350 $Y=110020 $dt=4
Q15 GNDA GNDA 21 qpvc3 $X=319350 $Y=126770 $dt=4
Q16 GNDA GNDA 21 qpvc3 $X=336105 $Y=9520 $dt=4
Q17 GNDA GNDA 21 qpvc3 $X=336105 $Y=26270 $dt=4
Q18 GNDA GNDA 21 qpvc3 $X=336105 $Y=43020 $dt=4
Q19 GNDA GNDA 21 qpvc3 $X=336105 $Y=59770 $dt=4
Q20 GNDA GNDA 21 qpvc3 $X=336105 $Y=76520 $dt=4
Q21 GNDA GNDA 21 qpvc3 $X=336105 $Y=93270 $dt=4
Q22 GNDA GNDA 21 qpvc3 $X=336105 $Y=110020 $dt=4
Q23 GNDA GNDA 21 qpvc3 $X=336105 $Y=126770 $dt=4
Q24 GNDA GNDA 21 qpvc3 $X=352860 $Y=9520 $dt=4
Q25 GNDA GNDA 21 qpvc3 $X=352860 $Y=26270 $dt=4
Q26 GNDA GNDA 21 qpvc3 $X=352860 $Y=43020 $dt=4
Q27 GNDA GNDA 21 qpvc3 $X=352860 $Y=59770 $dt=4
Q28 GNDA GNDA 21 qpvc3 $X=352860 $Y=76520 $dt=4
Q29 GNDA GNDA 21 qpvc3 $X=352860 $Y=93270 $dt=4
Q30 GNDA GNDA 21 qpvc3 $X=352860 $Y=110020 $dt=4
Q31 GNDA GNDA 21 qpvc3 $X=352860 $Y=126770 $dt=4
D32 GNDA VDD3A p_dnw AREA=1.07147e-09 PJ=0.0001732 perimeter=0.0001732 $X=3950 $Y=96990 $dt=5
D33 GNDA VDD3A p_dnw AREA=2.50005e-10 PJ=8.653e-05 perimeter=8.653e-05 $X=6985 $Y=72595 $dt=5
D34 GNDA VDD3A p_dnw AREA=1.35123e-09 PJ=0.00022788 perimeter=0.00022788 $X=35895 $Y=52775 $dt=5
D35 GNDA VDD3A p_dnw AREA=3.30547e-10 PJ=0.00010554 perimeter=0.00010554 $X=57005 $Y=102040 $dt=5
D36 GNDA VDD3A p_dnw AREA=1.64117e-10 PJ=7.372e-05 perimeter=7.372e-05 $X=76425 $Y=117950 $dt=5
D37 GNDA VDD3A p_dnw AREA=1.17512e-09 PJ=0.00013712 perimeter=0.00013712 $X=119255 $Y=7325 $dt=5
D38 GNDA VDD3A p_dnw3 AREA=3.99668e-10 PJ=0 perimeter=0 $X=9150 $Y=105110 $dt=8
D39 GNDA VDD3A p_dnw3 AREA=3.99668e-10 PJ=0 perimeter=0 $X=9150 $Y=118090 $dt=8
D40 GNDA VDD3A p_dnw3 AREA=7.74011e-10 PJ=0 perimeter=0 $X=41595 $Y=59115 $dt=8
D41 GNDA VDD3A p_dnw3 AREA=7.74011e-10 PJ=0 perimeter=0 $X=41595 $Y=72735 $dt=8
D42 GNDA VDD3A p_dnw3 AREA=1.71976e-10 PJ=0 perimeter=0 $X=58145 $Y=118370 $dt=8
D43 GNDA VDD3A p_dnw3 AREA=1.71976e-10 PJ=0 perimeter=0 $X=77565 $Y=124290 $dt=8
C44 14 OUT area=9e-10 perimeter=0.00012 $[cmm5t] $X=121395 $Y=9465 $dt=11
.ends bandgap_su

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: mosvc3_CDNS_7246542145921                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt mosvc3_CDNS_7246542145921 1 2
** N=2 EP=2 FDC=2
X0 2 1 1 MOSVC3 w=2.5e-05 l=3e-05 $X=0 $Y=0 $dt=3
D1 1 1 p_dnw3 AREA=6.7176e-11 PJ=0.00011492 perimeter=0.00011492 $X=-800 $Y=-430 $dt=8
.ends mosvc3_CDNS_7246542145921

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3i_6_CDNS_7246542145922                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3i_6_CDNS_7246542145922 1 2 3
** N=3 EP=3 FDC=4
X0 1 3 3 1 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=4.8e-12 ps=1.054e-05 pd=2.096e-05 $X=0 $Y=0 $dt=2
X1 3 3 1 1 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=4.8e-12 ad=2.7e-12 ps=2.096e-05 pd=1.054e-05 $X=3040 $Y=0 $dt=2
D2 1 2 p_ddnw AREA=3.07331e-10 PJ=7.576e-05 perimeter=7.576e-05 $X=-6110 $Y=-4940 $dt=6
D3 1 2 p_dipdnwmv AREA=7.49452e-11 PJ=4.496e-05 perimeter=4.496e-05 $X=-2260 $Y=-1090 $dt=7
.ends ne3i_6_CDNS_7246542145922

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246542145923                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246542145923 1 2 3
** N=3 EP=3 FDC=2
M0 2 2 1 1 pe3 L=1e-05 W=2e-06 AD=9.6e-13 AS=9.6e-13 PD=4.96e-06 PS=4.96e-06 $X=0 $Y=0 $dt=1
D1 3 1 p_dnw3 AREA=4.57434e-11 PJ=3.138e-05 perimeter=3.138e-05 $X=-910 $Y=-1440 $dt=8
.ends pe3_CDNS_7246542145923

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_7246542145924                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_7246542145924 1 2 3 4
** N=4 EP=4 FDC=2
M0 3 2 1 4 ne3 L=2.5e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
M1 1 2 3 4 ne3 L=2.5e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=3040 $Y=0 $dt=0
.ends ne3_CDNS_7246542145924

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246542145925                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246542145925 1 2 3 4 5
** N=5 EP=5 FDC=3
M0 3 2 1 4 pe3 L=2.5e-06 W=1e-05 AD=2.7e-12 AS=4.8e-12 PD=1.054e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
M1 1 2 3 4 pe3 L=2.5e-06 W=1e-05 AD=4.8e-12 AS=2.7e-12 PD=2.096e-05 PS=1.054e-05 $X=3040 $Y=0 $dt=1
D2 5 4 p_dnw3 AREA=1.03234e-10 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=8
.ends pe3_CDNS_7246542145925

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246542145926                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246542145926 1 2 3 4 5
** N=5 EP=5 FDC=2
M0 3 2 1 4 pe3 L=2.5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
D1 5 4 p_dnw3 AREA=6.65712e-11 PJ=0 perimeter=0 $X=-1510 $Y=-1030 $dt=8
.ends pe3_CDNS_7246542145926

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_7246542145927                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_7246542145927 1 2 3
*.DEVICECLIMB
** N=4 EP=3 FDC=1
M0 3 2 1 1 pe3 L=2.5e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_7246542145927

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3i_6_CDNS_7246542145928                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3i_6_CDNS_7246542145928 1 2 3 4 5
** N=5 EP=5 FDC=10
X0 3 4 5 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=4.8e-12 ps=1.054e-05 pd=2.096e-05 $X=0 $Y=0 $dt=2
X1 5 4 3 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=2.7e-12 ps=1.054e-05 pd=1.054e-05 $X=3040 $Y=0 $dt=2
X2 3 4 5 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=2.7e-12 ps=1.054e-05 pd=1.054e-05 $X=6080 $Y=0 $dt=2
X3 5 4 3 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=2.7e-12 ps=1.054e-05 pd=1.054e-05 $X=9120 $Y=0 $dt=2
X4 3 4 5 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=2.7e-12 ps=1.054e-05 pd=1.054e-05 $X=12160 $Y=0 $dt=2
X5 5 4 3 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=2.7e-12 ps=1.054e-05 pd=1.054e-05 $X=15200 $Y=0 $dt=2
X6 3 4 5 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=2.7e-12 ad=2.7e-12 ps=1.054e-05 pd=1.054e-05 $X=18240 $Y=0 $dt=2
X7 5 4 3 3 2 1 NE3I_6 w=1e-05 l=2.5e-06 as=4.8e-12 ad=2.7e-12 ps=2.096e-05 pd=1.054e-05 $X=21280 $Y=0 $dt=2
D8 1 2 p_ddnw AREA=5.2432e-10 PJ=0.00011224 perimeter=0.00011224 $X=-6110 $Y=-4940 $dt=6
D9 3 2 p_dipdnwmv AREA=1.51486e-10 PJ=8.144e-05 perimeter=8.144e-05 $X=-2260 $Y=-1090 $dt=7
.ends ne3i_6_CDNS_7246542145928

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_7246542145929                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_7246542145929 1 2 3
*.DEVICECLIMB
** N=3 EP=3 FDC=1
R0 2 1 L=0.0002878 W=4e-06 $[rpp1k1_3] $SUB=3 $X=-4220 $Y=0 $dt=10
.ends rpp1k1_3_CDNS_7246542145929

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: constant_gm                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt constant_gm GNDA VDD3 OUT1 OUT2 OUT3
** N=16 EP=5 FDC=56
X94 GNDA VDD3 13 ne3i_6_CDNS_7246542145922 $T=18020 14875 0 0 $X=7250 $Y=5275
X95 16 12 GNDA pe3_CDNS_7246542145923 $T=10155 41775 0 0 $X=8645 $Y=39735
X96 11 16 GNDA pe3_CDNS_7246542145923 $T=20155 47905 1 180 $X=8645 $Y=45865
X97 13 12 12 GNDA ne3_CDNS_7246542145924 $T=25460 39505 0 0 $X=24660 $Y=39105
X98 14 12 11 GNDA ne3_CDNS_7246542145924 $T=34790 39505 0 0 $X=33990 $Y=39105
X99 6 11 12 VDD3 GNDA pe3_CDNS_7246542145925 $T=11660 58745 0 0 $X=10150 $Y=57715
X100 7 11 11 VDD3 GNDA pe3_CDNS_7246542145925 $T=21810 58745 0 0 $X=20300 $Y=57715
X101 8 11 OUT1 VDD3 GNDA pe3_CDNS_7246542145925 $T=32565 58745 0 0 $X=31055 $Y=57715
X102 9 11 OUT2 VDD3 GNDA pe3_CDNS_7246542145925 $T=43380 58745 0 0 $X=41870 $Y=57715
X103 10 11 OUT3 VDD3 GNDA pe3_CDNS_7246542145926 $T=53845 58745 0 0 $X=52335 $Y=57715
X104 VDD3 VDD3 VDD3 pe3_CDNS_7246542145927 $T=18765 87600 1 0 $X=17255 $Y=76570
X105 VDD3 VDD3 VDD3 pe3_CDNS_7246542145927 $T=18765 106960 1 0 $X=17255 $Y=95930
X106 VDD3 7 9 pe3_CDNS_7246542145927 $T=22505 87600 1 0 $X=20995 $Y=76570
X107 VDD3 7 9 pe3_CDNS_7246542145927 $T=22505 106960 1 0 $X=20995 $Y=95930
X108 VDD3 7 7 pe3_CDNS_7246542145927 $T=26245 87600 1 0 $X=24735 $Y=76570
X109 VDD3 7 6 pe3_CDNS_7246542145927 $T=26245 106960 1 0 $X=24735 $Y=95930
X110 VDD3 7 6 pe3_CDNS_7246542145927 $T=29985 87600 1 0 $X=28475 $Y=76570
X111 VDD3 7 7 pe3_CDNS_7246542145927 $T=29985 106960 1 0 $X=28475 $Y=95930
X112 VDD3 7 8 pe3_CDNS_7246542145927 $T=33725 87600 1 0 $X=32215 $Y=76570
X113 VDD3 7 8 pe3_CDNS_7246542145927 $T=33725 106960 1 0 $X=32215 $Y=95930
X114 VDD3 VDD3 VDD3 pe3_CDNS_7246542145927 $T=37465 87600 1 0 $X=35955 $Y=76570
X115 VDD3 7 10 pe3_CDNS_7246542145927 $T=37465 106960 1 0 $X=35955 $Y=95930
X116 VDD3 VDD3 VDD3 pe3_CDNS_7246542145927 $T=41205 87600 1 0 $X=39695 $Y=76570
X117 VDD3 VDD3 VDD3 pe3_CDNS_7246542145927 $T=41205 106960 1 0 $X=39695 $Y=95930
X118 GNDA VDD3 15 13 14 ne3i_6_CDNS_7246542145928 $T=48275 14875 0 0 $X=37505 $Y=5275
X119 GNDA 15 VDD3 rpp1k1_3_CDNS_7246542145929 $T=62765 46455 1 90 $X=62545 $Y=41295
D0 GNDA VDD3 p_dnw AREA=4.77568e-10 PJ=0.00014131 perimeter=0.00014131 $X=7700 $Y=53605 $dt=5
D1 GNDA VDD3 p_dnw AREA=1.16854e-09 PJ=0.00017172 perimeter=0.00017172 $X=12555 $Y=74150 $dt=5
D2 GNDA VDD3 p_dnw AREA=1.48411e-09 PJ=0.00019385 perimeter=0.00019385 $X=61625 $Y=40375 $dt=5
D3 GNDA VDD3 p_dnw3 AREA=3.37198e-10 PJ=0 perimeter=0 $X=17255 $Y=76570 $dt=8
D4 GNDA VDD3 p_dnw3 AREA=3.37198e-10 PJ=0 perimeter=0 $X=17255 $Y=95930 $dt=8
.ends constant_gm

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: bias                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt bias BGAP_REF BIAS1 BIAS2 BIAS3 GNDA RES_BIAS VDDA
** N=9 EP=7 FDC=460
X1 GNDA VDDA 1 RES_BIAS BIAS2 BIAS1 BGAP_REF ref_bias $T=469540 4625 0 0 $X=471000 $Y=6590
X2 GNDA VDDA 8 BGAP_REF bandgap_su $T=97685 3355 0 0 $X=99220 $Y=6370
X3 GNDA VDDA mosvc3_CDNS_7246542145921 $T=25775 183420 1 0 $X=24975 $Y=157800
X4 GNDA VDDA mosvc3_CDNS_7246542145921 $T=25775 185680 0 0 $X=24975 $Y=185250
X5 GNDA VDDA mosvc3_CDNS_7246542145921 $T=58775 183420 1 0 $X=57975 $Y=157800
X6 GNDA VDDA mosvc3_CDNS_7246542145921 $T=58775 185680 0 0 $X=57975 $Y=185250
X7 GNDA VDDA mosvc3_CDNS_7246542145921 $T=91775 183420 1 0 $X=90975 $Y=157800
X8 GNDA VDDA mosvc3_CDNS_7246542145921 $T=91775 185680 0 0 $X=90975 $Y=185250
X9 GNDA VDDA mosvc3_CDNS_7246542145921 $T=124775 183420 1 0 $X=123975 $Y=157800
X10 GNDA VDDA mosvc3_CDNS_7246542145921 $T=124775 185680 0 0 $X=123975 $Y=185250
X11 GNDA VDDA mosvc3_CDNS_7246542145921 $T=157775 183420 1 0 $X=156975 $Y=157800
X12 GNDA VDDA mosvc3_CDNS_7246542145921 $T=157775 185680 0 0 $X=156975 $Y=185250
X13 GNDA VDDA mosvc3_CDNS_7246542145921 $T=190775 183420 1 0 $X=189975 $Y=157800
X14 GNDA VDDA mosvc3_CDNS_7246542145921 $T=190775 185680 0 0 $X=189975 $Y=185250
X15 GNDA VDDA mosvc3_CDNS_7246542145921 $T=223775 183420 1 0 $X=222975 $Y=157800
X16 GNDA VDDA mosvc3_CDNS_7246542145921 $T=223775 185680 0 0 $X=222975 $Y=185250
X17 GNDA VDDA mosvc3_CDNS_7246542145921 $T=256775 183420 1 0 $X=255975 $Y=157800
X18 GNDA VDDA mosvc3_CDNS_7246542145921 $T=256775 185680 0 0 $X=255975 $Y=185250
X19 GNDA VDDA mosvc3_CDNS_7246542145921 $T=289775 183420 1 0 $X=288975 $Y=157800
X20 GNDA VDDA mosvc3_CDNS_7246542145921 $T=289775 185680 0 0 $X=288975 $Y=185250
X21 GNDA VDDA mosvc3_CDNS_7246542145921 $T=322775 183420 1 0 $X=321975 $Y=157800
X22 GNDA VDDA mosvc3_CDNS_7246542145921 $T=322775 185680 0 0 $X=321975 $Y=185250
X23 GNDA VDDA mosvc3_CDNS_7246542145921 $T=355775 183420 1 0 $X=354975 $Y=157800
X24 GNDA VDDA mosvc3_CDNS_7246542145921 $T=355775 185680 0 0 $X=354975 $Y=185250
X25 GNDA VDDA mosvc3_CDNS_7246542145921 $T=388775 183420 1 0 $X=387975 $Y=157800
X26 GNDA VDDA mosvc3_CDNS_7246542145921 $T=388775 185680 0 0 $X=387975 $Y=185250
X27 GNDA VDDA mosvc3_CDNS_7246542145921 $T=421775 183420 1 0 $X=420975 $Y=157800
X28 GNDA VDDA mosvc3_CDNS_7246542145921 $T=421775 185680 0 0 $X=420975 $Y=185250
X29 GNDA VDDA 1 8 BIAS3 constant_gm $T=6360 5750 0 0 $X=7225 $Y=6590
.ends bias
