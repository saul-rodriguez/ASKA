* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : hvswitch8                                    *
* Netlisted  : Mon Aug 26 08:53:08 2024                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 LDDN(nedia) nedia2_d dnwtrm(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 1 LDDP(ped) ped12_d pwitrm(D) p1trm(G) pdiff(S) bulk(B)
*.DEVTMPLT 2 MN(ne3) nem ndiff(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 3 MP(pe3) pem pdiff(D) p1trm(G) pdiff(S) nwtrm(B)
*.DEVTMPLT 4 D(p_dnw) p_dnw bulk(POS) nwtrm(NEG)
*.DEVTMPLT 5 D(p_ddnw) p_ddnw bulk(POS) dnwtrm(NEG)
*.DEVTMPLT 6 D(p_dwhn) p_dwhn bulk(POS) hnw(NEG)
*.DEVTMPLT 7 D(dpp20) dpp20 pwitrm(POS) dnwtrm(NEG)
*.DEVTMPLT 8 D(dsba) d_dsba d_dsdf(POS) hnw(NEG) bulk(SUB)
*.DEVTMPLT 9 D(p_dnw3) p_dnwm bulk(POS) nwtrm(NEG)
*.DEVTMPLT 10 R(rpp1k1_3) rpp1k1_s p1trm(POS) p1trm(NEG) bulk(SUB)
*.DEVTMPLT 11 C(csf4a) d_csf4a m1atrm(POS) m1btrm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246551802815                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246551802815 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246551802815

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246551802833                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246551802833 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246551802833

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246551802834                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246551802834 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246551802834

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246551802842                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246551802842 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246551802842

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246551802846                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246551802846 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246551802846

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246551802847                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246551802847 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246551802847

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246551802848                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246551802848 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246551802848

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246551802850                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246551802850 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246551802850

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246551802851                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246551802851 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246551802851

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246551802854                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246551802854 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246551802854

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246551802855                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246551802855 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246551802855

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nedia_CDNS_724655180280                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nedia_CDNS_724655180280 1 2 3 4
** N=4 EP=4 FDC=12
X0 2 3 4 1 LDDN w=5e-05 l=1.25e-06 adio=6.71697e-10 pdio=3.30958e-05 extlay=1 $[nedia] $X=-680 $Y=-4850 $dt=0
X1 2 3 4 1 LDDN w=5e-05 l=1.25e-06 adio=6.71697e-10 pdio=3.30958e-05 extlay=1 $[nedia] $X=11220 $Y=-4850 $dt=0
X2 2 3 4 1 LDDN w=5e-05 l=1.25e-06 adio=6.71697e-10 pdio=3.30958e-05 extlay=1 $[nedia] $X=23120 $Y=-4850 $dt=0
X3 2 3 4 1 LDDN w=5e-05 l=1.25e-06 adio=6.71697e-10 pdio=3.30958e-05 extlay=1 $[nedia] $X=35020 $Y=-4850 $dt=0
X4 2 3 4 1 LDDN w=5e-05 l=1.25e-06 adio=6.71697e-10 pdio=3.30958e-05 extlay=1 $[nedia] $X=46920 $Y=-4850 $dt=0
X5 2 3 4 1 LDDN w=5e-05 l=1.25e-06 adio=6.71697e-10 pdio=3.30958e-05 extlay=1 $[nedia] $X=58820 $Y=-4850 $dt=0
X6 2 3 4 1 LDDN w=5e-05 l=1.25e-06 adio=6.71697e-10 pdio=3.30958e-05 extlay=1 $[nedia] $X=70720 $Y=-4850 $dt=0
X7 2 3 4 1 LDDN w=5e-05 l=1.25e-06 adio=6.71697e-10 pdio=3.30958e-05 extlay=1 $[nedia] $X=82620 $Y=-4850 $dt=0
X8 2 3 4 1 LDDN w=5e-05 l=1.25e-06 adio=6.71697e-10 pdio=3.30958e-05 extlay=1 $[nedia] $X=94520 $Y=-4850 $dt=0
X9 2 3 4 1 LDDN w=5e-05 l=1.25e-06 adio=6.71697e-10 pdio=3.30958e-05 extlay=1 $[nedia] $X=106420 $Y=-4850 $dt=0
X10 2 3 4 1 LDDN w=5e-05 l=1.25e-06 adio=6.71697e-10 pdio=3.30958e-05 extlay=1 $[nedia] $X=118320 $Y=-4850 $dt=0
X11 2 3 4 1 LDDN w=5e-05 l=1.25e-06 adio=6.71697e-10 pdio=3.30958e-05 extlay=1 $[nedia] $X=130220 $Y=-4850 $dt=0
.ends nedia_CDNS_724655180280

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X10                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X10 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7246551802815 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7246551802815 $T=500 1500 0 0 $X=0 $Y=1000
X2 1 VIATP_C_CDNS_7246551802815 $T=500 2500 0 0 $X=0 $Y=2000
X3 1 VIATP_C_CDNS_7246551802815 $T=500 3500 0 0 $X=0 $Y=3000
X4 1 VIATP_C_CDNS_7246551802815 $T=500 4500 0 0 $X=0 $Y=4000
X5 1 VIATP_C_CDNS_7246551802815 $T=500 5500 0 0 $X=0 $Y=5000
X6 1 VIATP_C_CDNS_7246551802815 $T=500 6500 0 0 $X=0 $Y=6000
X7 1 VIATP_C_CDNS_7246551802815 $T=500 7500 0 0 $X=0 $Y=7000
X8 1 VIATP_C_CDNS_7246551802815 $T=500 8500 0 0 $X=0 $Y=8000
X9 1 VIATP_C_CDNS_7246551802815 $T=500 9500 0 0 $X=0 $Y=9000
.ends MASCO__X10

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X12                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X12 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7246551802815 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7246551802815 $T=500 2500 0 0 $X=0 $Y=2000
X2 1 VIATP_C_CDNS_7246551802815 $T=500 4500 0 0 $X=0 $Y=4000
X3 1 VIATP_C_CDNS_7246551802815 $T=500 6500 0 0 $X=0 $Y=6000
X4 1 VIATP_C_CDNS_7246551802815 $T=500 8500 0 0 $X=0 $Y=8000
.ends MASCO__X12

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y19                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y19 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7246551802833 $T=500 620 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7246551802833 $T=1500 620 0 0 $X=1000 $Y=0
X2 1 VIATP_C_CDNS_7246551802833 $T=2500 620 0 0 $X=2000 $Y=0
X3 1 VIATP_C_CDNS_7246551802833 $T=3500 620 0 0 $X=3000 $Y=0
X4 1 VIATP_C_CDNS_7246551802833 $T=4500 620 0 0 $X=4000 $Y=0
X5 1 VIATP_C_CDNS_7246551802833 $T=5500 620 0 0 $X=5000 $Y=0
X6 1 VIATP_C_CDNS_7246551802833 $T=6500 620 0 0 $X=6000 $Y=0
X7 1 VIATP_C_CDNS_7246551802833 $T=7500 620 0 0 $X=7000 $Y=0
X8 1 VIATP_C_CDNS_7246551802833 $T=8500 620 0 0 $X=8000 $Y=0
X9 1 VIATP_C_CDNS_7246551802833 $T=9500 620 0 0 $X=9000 $Y=0
X10 1 VIATP_C_CDNS_7246551802833 $T=10500 620 0 0 $X=10000 $Y=0
X11 1 VIATP_C_CDNS_7246551802833 $T=11500 620 0 0 $X=11000 $Y=0
.ends MASCO__Y19

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y23                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y23 1
** N=1 EP=1 FDC=0
X0 1 MASCO__X12 $T=0 0 0 0 $X=0 $Y=0
X1 1 MASCO__X12 $T=2000 0 0 0 $X=2000 $Y=0
X2 1 MASCO__X12 $T=4000 0 0 0 $X=4000 $Y=0
X3 1 MASCO__X12 $T=6000 0 0 0 $X=6000 $Y=0
X4 1 MASCO__X12 $T=8000 0 0 0 $X=8000 $Y=0
X5 1 MASCO__X12 $T=10000 0 0 0 $X=10000 $Y=0
X6 1 MASCO__X12 $T=12000 0 0 0 $X=12000 $Y=0
X7 1 MASCO__X12 $T=14000 0 0 0 $X=14000 $Y=0
.ends MASCO__Y23

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y24                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y24 1
** N=1 EP=1 FDC=0
X0 1 MASCO__X10 $T=0 0 0 0 $X=0 $Y=0
X1 1 MASCO__X10 $T=2000 0 0 0 $X=2000 $Y=0
X2 1 MASCO__X10 $T=4000 0 0 0 $X=4000 $Y=0
X3 1 MASCO__X10 $T=6000 0 0 0 $X=6000 $Y=0
X4 1 MASCO__X10 $T=8000 0 0 0 $X=8000 $Y=0
X5 1 MASCO__X10 $T=10000 0 0 0 $X=10000 $Y=0
X6 1 MASCO__X10 $T=12000 0 0 0 $X=12000 $Y=0
X7 1 MASCO__X10 $T=14000 0 0 0 $X=14000 $Y=0
.ends MASCO__Y24

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__H1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__H1 1 2 3 4
** N=4 EP=4 FDC=12
X0 4 VIATP_C_CDNS_7246551802815 $T=346380 92210 0 0 $X=345880 $Y=91710
X1 4 VIATP_C_CDNS_7246551802833 $T=234380 102330 0 0 $X=233880 $Y=101710
X2 3 VIATP_C_CDNS_7246551802833 $T=257995 144490 0 0 $X=257495 $Y=143870
X3 3 VIATP_C_CDNS_7246551802833 $T=258995 144490 0 0 $X=258495 $Y=143870
X4 3 VIATP_C_CDNS_7246551802833 $T=259995 144490 0 0 $X=259495 $Y=143870
X5 3 VIATP_C_CDNS_7246551802833 $T=260995 144490 0 0 $X=260495 $Y=143870
X6 3 VIATP_C_CDNS_7246551802833 $T=261995 144490 0 0 $X=261495 $Y=143870
X7 3 VIATP_C_CDNS_7246551802833 $T=262995 144490 0 0 $X=262495 $Y=143870
X8 3 VIATP_C_CDNS_7246551802833 $T=263995 144490 0 0 $X=263495 $Y=143870
X9 3 VIATP_C_CDNS_7246551802833 $T=264995 144490 0 0 $X=264495 $Y=143870
X10 3 VIATP_C_CDNS_7246551802833 $T=265995 144490 0 0 $X=265495 $Y=143870
X11 3 VIATP_C_CDNS_7246551802833 $T=266995 144490 0 0 $X=266495 $Y=143870
X12 4 VIATP_C_CDNS_7246551802833 $T=343380 102330 0 0 $X=342880 $Y=101710
X13 4 VIATP_C_CDNS_7246551802833 $T=344380 102330 0 0 $X=343880 $Y=101710
X14 4 VIATP_C_CDNS_7246551802833 $T=345380 102330 0 0 $X=344880 $Y=101710
X15 3 VIATP_C_CDNS_7246551802833 $T=365995 144490 0 0 $X=365495 $Y=143870
X16 3 VIATP_C_CDNS_7246551802833 $T=366995 144490 0 0 $X=366495 $Y=143870
X17 3 VIATP_C_CDNS_7246551802833 $T=367995 144490 0 0 $X=367495 $Y=143870
X18 3 VIATP_C_CDNS_7246551802833 $T=368995 144490 0 0 $X=368495 $Y=143870
X19 3 VIATP_C_CDNS_7246551802833 $T=369995 144490 0 0 $X=369495 $Y=143870
X20 3 VIATP_C_CDNS_7246551802833 $T=370995 144490 0 0 $X=370495 $Y=143870
X21 3 VIATP_C_CDNS_7246551802833 $T=371995 144490 0 0 $X=371495 $Y=143870
X22 4 VIATP_C_CDNS_7246551802833 $T=372380 102330 0 0 $X=371880 $Y=101710
X23 3 VIATP_C_CDNS_7246551802833 $T=372995 144490 0 0 $X=372495 $Y=143870
X24 4 VIATP_C_CDNS_7246551802833 $T=373380 102330 0 0 $X=372880 $Y=101710
X25 3 VIATP_C_CDNS_7246551802833 $T=373995 144490 0 0 $X=373495 $Y=143870
X26 4 VIATP_C_CDNS_7246551802833 $T=374380 102330 0 0 $X=373880 $Y=101710
X27 3 VIATP_C_CDNS_7246551802833 $T=374995 144490 0 0 $X=374495 $Y=143870
X28 4 VIATP_C_CDNS_7246551802833 $T=375380 102330 0 0 $X=374880 $Y=101710
X29 3 VIATP_C_CDNS_7246551802833 $T=375995 144490 0 0 $X=375495 $Y=143870
X30 4 VIATP_C_CDNS_7246551802833 $T=376380 102330 0 0 $X=375880 $Y=101710
X31 3 VIATP_C_CDNS_7246551802833 $T=377995 144490 0 0 $X=377495 $Y=143870
X32 4 VIATP_C_CDNS_7246551802833 $T=378380 102330 0 0 $X=377880 $Y=101710
X33 3 VIATP_C_CDNS_7246551802833 $T=378995 144490 0 0 $X=378495 $Y=143870
X34 4 VIATP_C_CDNS_7246551802833 $T=379380 102330 0 0 $X=378880 $Y=101710
X35 3 VIATP_C_CDNS_7246551802833 $T=379995 144490 0 0 $X=379495 $Y=143870
X36 4 VIATP_C_CDNS_7246551802833 $T=380380 102330 0 0 $X=379880 $Y=101710
X37 3 VIATP_C_CDNS_7246551802833 $T=380995 144490 0 0 $X=380495 $Y=143870
X38 4 VIATP_C_CDNS_7246551802833 $T=381380 102330 0 0 $X=380880 $Y=101710
X39 3 VIATP_C_CDNS_7246551802833 $T=381995 144490 0 0 $X=381495 $Y=143870
X40 4 VIATP_C_CDNS_7246551802833 $T=382380 102330 0 0 $X=381880 $Y=101710
X41 3 VIATP_C_CDNS_7246551802833 $T=382995 144490 0 0 $X=382495 $Y=143870
X42 4 VIATP_C_CDNS_7246551802833 $T=383380 102330 0 0 $X=382880 $Y=101710
X43 3 VIATP_C_CDNS_7246551802833 $T=383995 144490 0 0 $X=383495 $Y=143870
X44 4 VIATP_C_CDNS_7246551802833 $T=384380 102330 0 0 $X=383880 $Y=101710
X45 3 VIATP_C_CDNS_7246551802833 $T=384995 144490 0 0 $X=384495 $Y=143870
X46 4 VIATP_C_CDNS_7246551802833 $T=385380 102330 0 0 $X=384880 $Y=101710
X47 4 VIATP_C_CDNS_7246551802834 $T=377440 102330 0 0 $X=377000 $Y=101710
X48 3 VIATP_C_CDNS_7246551802842 $T=376745 145610 0 0 $X=376475 $Y=145110
X49 3 VIATP_C_CDNS_7246551802842 $T=376745 146610 0 0 $X=376475 $Y=146110
X50 3 VIATP_C_CDNS_7246551802842 $T=376745 147610 0 0 $X=376475 $Y=147110
X51 3 VIATP_C_CDNS_7246551802842 $T=376745 148610 0 0 $X=376475 $Y=148110
X52 3 VIATP_C_CDNS_7246551802842 $T=376745 149610 0 0 $X=376475 $Y=149110
X53 3 VIATP_C_CDNS_7246551802842 $T=376745 150610 0 0 $X=376475 $Y=150110
X54 3 VIATP_C_CDNS_7246551802842 $T=376745 151610 0 0 $X=376475 $Y=151110
X55 3 VIATP_C_CDNS_7246551802842 $T=376745 152610 0 0 $X=376475 $Y=152110
X56 3 VIATP_C_CDNS_7246551802842 $T=376745 153610 0 0 $X=376475 $Y=153110
X57 3 VIATP_C_CDNS_7246551802842 $T=376745 154610 0 0 $X=376475 $Y=154110
X58 3 VIATP_C_CDNS_7246551802846 $T=232755 144490 0 0 $X=232025 $Y=143870
X59 3 VIATP_C_CDNS_7246551802847 $T=268645 145610 0 0 $X=268375 $Y=145110
X60 3 VIATP_C_CDNS_7246551802847 $T=268645 146610 0 0 $X=268375 $Y=146110
X61 3 VIATP_C_CDNS_7246551802847 $T=268645 147610 0 0 $X=268375 $Y=147110
X62 3 VIATP_C_CDNS_7246551802847 $T=268645 148610 0 0 $X=268375 $Y=148110
X63 3 VIATP_C_CDNS_7246551802847 $T=268645 149610 0 0 $X=268375 $Y=149110
X64 3 VIATP_C_CDNS_7246551802847 $T=268645 150610 0 0 $X=268375 $Y=150110
X65 3 VIATP_C_CDNS_7246551802847 $T=268645 151610 0 0 $X=268375 $Y=151110
X66 3 VIATP_C_CDNS_7246551802847 $T=268645 152610 0 0 $X=268375 $Y=152110
X67 3 VIATP_C_CDNS_7246551802847 $T=268645 153610 0 0 $X=268375 $Y=153110
X68 3 VIATP_C_CDNS_7246551802847 $T=268645 154610 0 0 $X=268375 $Y=154110
X69 3 VIATP_C_CDNS_7246551802848 $T=232755 145610 0 0 $X=232025 $Y=145110
X70 3 VIATP_C_CDNS_7246551802848 $T=232755 146610 0 0 $X=232025 $Y=146110
X71 3 VIATP_C_CDNS_7246551802848 $T=232755 147610 0 0 $X=232025 $Y=147110
X72 3 VIATP_C_CDNS_7246551802848 $T=232755 148610 0 0 $X=232025 $Y=148110
X73 3 VIATP_C_CDNS_7246551802848 $T=232755 149610 0 0 $X=232025 $Y=149110
X74 3 VIATP_C_CDNS_7246551802848 $T=232755 150610 0 0 $X=232025 $Y=150110
X75 3 VIATP_C_CDNS_7246551802848 $T=232755 151610 0 0 $X=232025 $Y=151110
X76 3 VIATP_C_CDNS_7246551802848 $T=232755 152610 0 0 $X=232025 $Y=152110
X77 3 VIATP_C_CDNS_7246551802848 $T=232755 153610 0 0 $X=232025 $Y=153110
X78 3 VIATP_C_CDNS_7246551802848 $T=232755 154610 0 0 $X=232025 $Y=154110
X79 4 VIATP_C_CDNS_7246551802850 $T=232950 102330 0 0 $X=232020 $Y=101710
X80 4 VIATP_C_CDNS_7246551802851 $T=232950 92210 0 0 $X=232020 $Y=91710
X81 4 VIATP_C_CDNS_7246551802851 $T=232950 93210 0 0 $X=232020 $Y=92710
X82 4 VIATP_C_CDNS_7246551802851 $T=232950 94210 0 0 $X=232020 $Y=93710
X83 4 VIATP_C_CDNS_7246551802851 $T=232950 95210 0 0 $X=232020 $Y=94710
X84 4 VIATP_C_CDNS_7246551802851 $T=232950 96210 0 0 $X=232020 $Y=95710
X85 4 VIATP_C_CDNS_7246551802851 $T=232950 97210 0 0 $X=232020 $Y=96710
X86 4 VIATP_C_CDNS_7246551802851 $T=232950 98210 0 0 $X=232020 $Y=97710
X87 4 VIATP_C_CDNS_7246551802851 $T=232950 99210 0 0 $X=232020 $Y=98710
X88 4 VIATP_C_CDNS_7246551802851 $T=232950 100210 0 0 $X=232020 $Y=99710
X89 4 VIATP_C_CDNS_7246551802851 $T=232950 101210 0 0 $X=232020 $Y=100710
X90 4 VIATP_C_CDNS_7246551802854 $T=377440 92210 0 0 $X=377000 $Y=91710
X91 4 VIATP_C_CDNS_7246551802854 $T=377440 93210 0 0 $X=377000 $Y=92710
X92 4 VIATP_C_CDNS_7246551802854 $T=377440 94210 0 0 $X=377000 $Y=93710
X93 4 VIATP_C_CDNS_7246551802854 $T=377440 95210 0 0 $X=377000 $Y=94710
X94 4 VIATP_C_CDNS_7246551802854 $T=377440 96210 0 0 $X=377000 $Y=95710
X95 4 VIATP_C_CDNS_7246551802854 $T=377440 97210 0 0 $X=377000 $Y=96710
X96 4 VIATP_C_CDNS_7246551802854 $T=377440 98210 0 0 $X=377000 $Y=97710
X97 4 VIATP_C_CDNS_7246551802854 $T=377440 99210 0 0 $X=377000 $Y=98710
X98 4 VIATP_C_CDNS_7246551802854 $T=377440 100210 0 0 $X=377000 $Y=99710
X99 4 VIATP_C_CDNS_7246551802854 $T=377440 101210 0 0 $X=377000 $Y=100710
X100 4 VIATP_C_CDNS_7246551802855 $T=346510 94210 0 0 $X=346145 $Y=93710
X101 4 VIATP_C_CDNS_7246551802855 $T=346510 96210 0 0 $X=346145 $Y=95710
X102 4 VIATP_C_CDNS_7246551802855 $T=346510 98210 0 0 $X=346145 $Y=97710
X103 4 VIATP_C_CDNS_7246551802855 $T=346510 100210 0 0 $X=346145 $Y=99710
X104 1 3 2 4 nedia_CDNS_724655180280 $T=238930 110910 0 0 $X=222710 $Y=91520
X105 3 MASCO__X10 $T=234495 145110 0 0 $X=234495 $Y=145110
X106 3 MASCO__X10 $T=236495 145110 0 0 $X=236495 $Y=145110
X107 3 MASCO__X10 $T=238495 145110 0 0 $X=238495 $Y=145110
X108 3 MASCO__X10 $T=240495 145110 0 0 $X=240495 $Y=145110
X109 3 MASCO__X10 $T=242495 145110 0 0 $X=242495 $Y=145110
X110 3 MASCO__X10 $T=244495 145110 0 0 $X=244495 $Y=145110
X111 3 MASCO__X10 $T=246495 145110 0 0 $X=246495 $Y=145110
X112 3 MASCO__X10 $T=248495 145110 0 0 $X=248495 $Y=145110
X113 3 MASCO__X10 $T=250495 145110 0 0 $X=250495 $Y=145110
X114 3 MASCO__X10 $T=270495 145110 0 0 $X=270495 $Y=145110
X115 3 MASCO__X10 $T=272495 145110 0 0 $X=272495 $Y=145110
X116 3 MASCO__X10 $T=274495 145110 0 0 $X=274495 $Y=145110
X117 3 MASCO__X10 $T=276495 145110 0 0 $X=276495 $Y=145110
X118 3 MASCO__X10 $T=278495 145110 0 0 $X=278495 $Y=145110
X119 3 MASCO__X10 $T=280495 145110 0 0 $X=280495 $Y=145110
X120 3 MASCO__X10 $T=282495 145110 0 0 $X=282495 $Y=145110
X121 3 MASCO__X10 $T=284495 145110 0 0 $X=284495 $Y=145110
X122 3 MASCO__X10 $T=286495 145110 0 0 $X=286495 $Y=145110
X123 3 MASCO__X10 $T=288495 145110 0 0 $X=288495 $Y=145110
X124 3 MASCO__X10 $T=290495 145110 0 0 $X=290495 $Y=145110
X125 3 MASCO__X10 $T=292495 145110 0 0 $X=292495 $Y=145110
X126 3 MASCO__X10 $T=294495 145110 0 0 $X=294495 $Y=145110
X127 3 MASCO__X10 $T=296495 145110 0 0 $X=296495 $Y=145110
X128 3 MASCO__X10 $T=298495 145110 0 0 $X=298495 $Y=145110
X129 3 MASCO__X10 $T=300495 145110 0 0 $X=300495 $Y=145110
X130 3 MASCO__X10 $T=302495 145110 0 0 $X=302495 $Y=145110
X131 3 MASCO__X10 $T=304495 145110 0 0 $X=304495 $Y=145110
X132 3 MASCO__X10 $T=306495 145110 0 0 $X=306495 $Y=145110
X133 3 MASCO__X10 $T=308495 145110 0 0 $X=308495 $Y=145110
X134 3 MASCO__X10 $T=310495 145110 0 0 $X=310495 $Y=145110
X135 3 MASCO__X10 $T=312495 145110 0 0 $X=312495 $Y=145110
X136 3 MASCO__X10 $T=314495 145110 0 0 $X=314495 $Y=145110
X137 3 MASCO__X10 $T=316495 145110 0 0 $X=316495 $Y=145110
X138 3 MASCO__X10 $T=318495 145110 0 0 $X=318495 $Y=145110
X139 3 MASCO__X10 $T=320495 145110 0 0 $X=320495 $Y=145110
X140 3 MASCO__X10 $T=322495 145110 0 0 $X=322495 $Y=145110
X141 3 MASCO__X10 $T=324495 145110 0 0 $X=324495 $Y=145110
X142 3 MASCO__X10 $T=326495 145110 0 0 $X=326495 $Y=145110
X143 3 MASCO__X10 $T=328495 145110 0 0 $X=328495 $Y=145110
X144 3 MASCO__X10 $T=330495 145110 0 0 $X=330495 $Y=145110
X145 3 MASCO__X10 $T=332495 145110 0 0 $X=332495 $Y=145110
X146 3 MASCO__X10 $T=334495 145110 0 0 $X=334495 $Y=145110
X147 3 MASCO__X10 $T=336495 145110 0 0 $X=336495 $Y=145110
X148 3 MASCO__X10 $T=338495 145110 0 0 $X=338495 $Y=145110
X149 3 MASCO__X10 $T=340495 145110 0 0 $X=340495 $Y=145110
X150 3 MASCO__X10 $T=342495 145110 0 0 $X=342495 $Y=145110
X151 3 MASCO__X10 $T=344495 145110 0 0 $X=344495 $Y=145110
X152 3 MASCO__X10 $T=346495 145110 0 0 $X=346495 $Y=145110
X153 3 MASCO__X10 $T=348495 145110 0 0 $X=348495 $Y=145110
X154 4 MASCO__X10 $T=348880 91710 0 0 $X=348880 $Y=91710
X155 3 MASCO__X10 $T=350495 145110 0 0 $X=350495 $Y=145110
X156 4 MASCO__X10 $T=350880 91710 0 0 $X=350880 $Y=91710
X157 3 MASCO__X10 $T=352495 145110 0 0 $X=352495 $Y=145110
X158 4 MASCO__X10 $T=352880 91710 0 0 $X=352880 $Y=91710
X159 3 MASCO__X10 $T=354495 145110 0 0 $X=354495 $Y=145110
X160 4 MASCO__X10 $T=354880 91710 0 0 $X=354880 $Y=91710
X161 3 MASCO__X10 $T=356495 145110 0 0 $X=356495 $Y=145110
X162 4 MASCO__X10 $T=356880 91710 0 0 $X=356880 $Y=91710
X163 3 MASCO__X10 $T=358495 145110 0 0 $X=358495 $Y=145110
X164 4 MASCO__X10 $T=358880 91710 0 0 $X=358880 $Y=91710
X165 3 MASCO__X10 $T=360495 145110 0 0 $X=360495 $Y=145110
X166 4 MASCO__X10 $T=360880 91710 0 0 $X=360880 $Y=91710
X167 3 MASCO__X10 $T=362495 145110 0 0 $X=362495 $Y=145110
X168 4 MASCO__X10 $T=362880 91710 0 0 $X=362880 $Y=91710
X169 3 MASCO__X10 $T=364495 145110 0 0 $X=364495 $Y=145110
X170 4 MASCO__X10 $T=364880 91710 0 0 $X=364880 $Y=91710
X171 3 MASCO__X10 $T=366495 145110 0 0 $X=366495 $Y=145110
X172 4 MASCO__X10 $T=366880 91710 0 0 $X=366880 $Y=91710
X173 3 MASCO__X10 $T=368495 145110 0 0 $X=368495 $Y=145110
X174 4 MASCO__X10 $T=368880 91710 0 0 $X=368880 $Y=91710
X175 3 MASCO__X10 $T=370495 145110 0 0 $X=370495 $Y=145110
X176 4 MASCO__X10 $T=370880 91710 0 0 $X=370880 $Y=91710
X177 3 MASCO__X10 $T=372495 145110 0 0 $X=372495 $Y=145110
X178 4 MASCO__X10 $T=372880 91710 0 0 $X=372880 $Y=91710
X179 3 MASCO__X10 $T=374495 145110 0 0 $X=374495 $Y=145110
X180 4 MASCO__X10 $T=374880 91710 0 0 $X=374880 $Y=91710
X181 3 MASCO__X10 $T=378495 145110 0 0 $X=378495 $Y=145110
X182 4 MASCO__X10 $T=378880 91710 0 0 $X=378880 $Y=91710
X183 3 MASCO__X10 $T=380495 145110 0 0 $X=380495 $Y=145110
X184 4 MASCO__X10 $T=380880 91710 0 0 $X=380880 $Y=91710
X185 3 MASCO__X10 $T=382495 145110 0 0 $X=382495 $Y=145110
X186 4 MASCO__X10 $T=382880 91710 0 0 $X=382880 $Y=91710
X187 3 MASCO__X10 $T=384495 145110 0 0 $X=384495 $Y=145110
X188 4 MASCO__X10 $T=384880 91710 0 0 $X=384880 $Y=91710
X189 3 MASCO__X12 $T=233495 146110 0 0 $X=233495 $Y=146110
X190 3 MASCO__X12 $T=235495 146110 0 0 $X=235495 $Y=146110
X191 3 MASCO__X12 $T=237495 146110 0 0 $X=237495 $Y=146110
X192 3 MASCO__X12 $T=239495 146110 0 0 $X=239495 $Y=146110
X193 3 MASCO__X12 $T=241495 146110 0 0 $X=241495 $Y=146110
X194 3 MASCO__X12 $T=243495 146110 0 0 $X=243495 $Y=146110
X195 3 MASCO__X12 $T=245495 146110 0 0 $X=245495 $Y=146110
X196 3 MASCO__X12 $T=247495 146110 0 0 $X=247495 $Y=146110
X197 3 MASCO__X12 $T=249495 146110 0 0 $X=249495 $Y=146110
X198 3 MASCO__X12 $T=269495 146110 0 0 $X=269495 $Y=146110
X199 3 MASCO__X12 $T=271495 146110 0 0 $X=271495 $Y=146110
X200 3 MASCO__X12 $T=273495 146110 0 0 $X=273495 $Y=146110
X201 3 MASCO__X12 $T=275495 146110 0 0 $X=275495 $Y=146110
X202 3 MASCO__X12 $T=277495 146110 0 0 $X=277495 $Y=146110
X203 3 MASCO__X12 $T=279495 146110 0 0 $X=279495 $Y=146110
X204 3 MASCO__X12 $T=281495 146110 0 0 $X=281495 $Y=146110
X205 3 MASCO__X12 $T=283495 146110 0 0 $X=283495 $Y=146110
X206 3 MASCO__X12 $T=285495 146110 0 0 $X=285495 $Y=146110
X207 3 MASCO__X12 $T=287495 146110 0 0 $X=287495 $Y=146110
X208 3 MASCO__X12 $T=289495 146110 0 0 $X=289495 $Y=146110
X209 3 MASCO__X12 $T=291495 146110 0 0 $X=291495 $Y=146110
X210 3 MASCO__X12 $T=293495 146110 0 0 $X=293495 $Y=146110
X211 3 MASCO__X12 $T=295495 146110 0 0 $X=295495 $Y=146110
X212 3 MASCO__X12 $T=297495 146110 0 0 $X=297495 $Y=146110
X213 3 MASCO__X12 $T=299495 146110 0 0 $X=299495 $Y=146110
X214 3 MASCO__X12 $T=301495 146110 0 0 $X=301495 $Y=146110
X215 3 MASCO__X12 $T=303495 146110 0 0 $X=303495 $Y=146110
X216 3 MASCO__X12 $T=305495 146110 0 0 $X=305495 $Y=146110
X217 3 MASCO__X12 $T=307495 146110 0 0 $X=307495 $Y=146110
X218 3 MASCO__X12 $T=309495 146110 0 0 $X=309495 $Y=146110
X219 3 MASCO__X12 $T=311495 146110 0 0 $X=311495 $Y=146110
X220 3 MASCO__X12 $T=313495 146110 0 0 $X=313495 $Y=146110
X221 3 MASCO__X12 $T=315495 146110 0 0 $X=315495 $Y=146110
X222 3 MASCO__X12 $T=317495 146110 0 0 $X=317495 $Y=146110
X223 3 MASCO__X12 $T=319495 146110 0 0 $X=319495 $Y=146110
X224 3 MASCO__X12 $T=321495 146110 0 0 $X=321495 $Y=146110
X225 3 MASCO__X12 $T=323495 146110 0 0 $X=323495 $Y=146110
X226 3 MASCO__X12 $T=325495 146110 0 0 $X=325495 $Y=146110
X227 3 MASCO__X12 $T=327495 146110 0 0 $X=327495 $Y=146110
X228 3 MASCO__X12 $T=329495 146110 0 0 $X=329495 $Y=146110
X229 3 MASCO__X12 $T=331495 146110 0 0 $X=331495 $Y=146110
X230 3 MASCO__X12 $T=333495 146110 0 0 $X=333495 $Y=146110
X231 3 MASCO__X12 $T=335495 146110 0 0 $X=335495 $Y=146110
X232 3 MASCO__X12 $T=337495 146110 0 0 $X=337495 $Y=146110
X233 3 MASCO__X12 $T=339495 146110 0 0 $X=339495 $Y=146110
X234 3 MASCO__X12 $T=341495 146110 0 0 $X=341495 $Y=146110
X235 3 MASCO__X12 $T=343495 146110 0 0 $X=343495 $Y=146110
X236 3 MASCO__X12 $T=345495 146110 0 0 $X=345495 $Y=146110
X237 3 MASCO__X12 $T=347495 146110 0 0 $X=347495 $Y=146110
X238 4 MASCO__X12 $T=347880 91710 0 0 $X=347880 $Y=91710
X239 3 MASCO__X12 $T=349495 146110 0 0 $X=349495 $Y=146110
X240 4 MASCO__X12 $T=349880 91710 0 0 $X=349880 $Y=91710
X241 3 MASCO__X12 $T=351495 146110 0 0 $X=351495 $Y=146110
X242 4 MASCO__X12 $T=351880 91710 0 0 $X=351880 $Y=91710
X243 3 MASCO__X12 $T=353495 146110 0 0 $X=353495 $Y=146110
X244 4 MASCO__X12 $T=353880 91710 0 0 $X=353880 $Y=91710
X245 3 MASCO__X12 $T=355495 146110 0 0 $X=355495 $Y=146110
X246 4 MASCO__X12 $T=355880 91710 0 0 $X=355880 $Y=91710
X247 3 MASCO__X12 $T=357495 146110 0 0 $X=357495 $Y=146110
X248 4 MASCO__X12 $T=357880 91710 0 0 $X=357880 $Y=91710
X249 3 MASCO__X12 $T=359495 146110 0 0 $X=359495 $Y=146110
X250 4 MASCO__X12 $T=359880 91710 0 0 $X=359880 $Y=91710
X251 3 MASCO__X12 $T=361495 146110 0 0 $X=361495 $Y=146110
X252 4 MASCO__X12 $T=361880 91710 0 0 $X=361880 $Y=91710
X253 3 MASCO__X12 $T=363495 146110 0 0 $X=363495 $Y=146110
X254 4 MASCO__X12 $T=363880 91710 0 0 $X=363880 $Y=91710
X255 3 MASCO__X12 $T=365495 146110 0 0 $X=365495 $Y=146110
X256 4 MASCO__X12 $T=365880 91710 0 0 $X=365880 $Y=91710
X257 3 MASCO__X12 $T=367495 146110 0 0 $X=367495 $Y=146110
X258 4 MASCO__X12 $T=367880 91710 0 0 $X=367880 $Y=91710
X259 3 MASCO__X12 $T=369495 146110 0 0 $X=369495 $Y=146110
X260 4 MASCO__X12 $T=369880 91710 0 0 $X=369880 $Y=91710
X261 3 MASCO__X12 $T=371495 146110 0 0 $X=371495 $Y=146110
X262 4 MASCO__X12 $T=371880 91710 0 0 $X=371880 $Y=91710
X263 3 MASCO__X12 $T=373495 146110 0 0 $X=373495 $Y=146110
X264 4 MASCO__X12 $T=373880 91710 0 0 $X=373880 $Y=91710
X265 4 MASCO__X12 $T=375880 91710 0 0 $X=375880 $Y=91710
X266 3 MASCO__X12 $T=377495 146110 0 0 $X=377495 $Y=146110
X267 4 MASCO__X12 $T=377880 91710 0 0 $X=377880 $Y=91710
X268 3 MASCO__X12 $T=379495 146110 0 0 $X=379495 $Y=146110
X269 4 MASCO__X12 $T=379880 91710 0 0 $X=379880 $Y=91710
X270 3 MASCO__X12 $T=381495 146110 0 0 $X=381495 $Y=146110
X271 4 MASCO__X12 $T=381880 91710 0 0 $X=381880 $Y=91710
X272 3 MASCO__X12 $T=383495 146110 0 0 $X=383495 $Y=146110
X273 4 MASCO__X12 $T=383880 91710 0 0 $X=383880 $Y=91710
X274 3 MASCO__Y19 $T=233495 143870 0 0 $X=233495 $Y=143870
X275 4 MASCO__Y19 $T=234880 101710 0 0 $X=234880 $Y=101710
X276 3 MASCO__Y19 $T=245495 143870 0 0 $X=245495 $Y=143870
X277 4 MASCO__Y19 $T=246880 101710 0 0 $X=246880 $Y=101710
X278 4 MASCO__Y19 $T=258880 101710 0 0 $X=258880 $Y=101710
X279 3 MASCO__Y19 $T=269495 143870 0 0 $X=269495 $Y=143870
X280 4 MASCO__Y19 $T=270880 101710 0 0 $X=270880 $Y=101710
X281 3 MASCO__Y19 $T=281495 143870 0 0 $X=281495 $Y=143870
X282 4 MASCO__Y19 $T=282880 101710 0 0 $X=282880 $Y=101710
X283 3 MASCO__Y19 $T=293495 143870 0 0 $X=293495 $Y=143870
X284 4 MASCO__Y19 $T=294880 101710 0 0 $X=294880 $Y=101710
X285 3 MASCO__Y19 $T=305495 143870 0 0 $X=305495 $Y=143870
X286 4 MASCO__Y19 $T=306880 101710 0 0 $X=306880 $Y=101710
X287 3 MASCO__Y19 $T=317495 143870 0 0 $X=317495 $Y=143870
X288 4 MASCO__Y19 $T=318880 101710 0 0 $X=318880 $Y=101710
X289 3 MASCO__Y19 $T=329495 143870 0 0 $X=329495 $Y=143870
X290 4 MASCO__Y19 $T=330880 101710 0 0 $X=330880 $Y=101710
X291 3 MASCO__Y19 $T=341495 143870 0 0 $X=341495 $Y=143870
X292 4 MASCO__Y19 $T=347880 101710 0 0 $X=347880 $Y=101710
X293 3 MASCO__Y19 $T=353495 143870 0 0 $X=353495 $Y=143870
X294 4 MASCO__Y19 $T=359880 101710 0 0 $X=359880 $Y=101710
X295 4 MASCO__Y23 $T=233880 91710 0 0 $X=233880 $Y=91710
X296 4 MASCO__Y23 $T=249880 91710 0 0 $X=249880 $Y=91710
X297 3 MASCO__Y23 $T=251495 146110 0 0 $X=251495 $Y=146110
X298 4 MASCO__Y23 $T=265880 91710 0 0 $X=265880 $Y=91710
X299 4 MASCO__Y23 $T=281880 91710 0 0 $X=281880 $Y=91710
X300 4 MASCO__Y23 $T=297880 91710 0 0 $X=297880 $Y=91710
X301 4 MASCO__Y23 $T=313880 91710 0 0 $X=313880 $Y=91710
X302 4 MASCO__Y23 $T=329880 91710 0 0 $X=329880 $Y=91710
X303 4 MASCO__Y24 $T=234880 91710 0 0 $X=234880 $Y=91710
X304 4 MASCO__Y24 $T=250880 91710 0 0 $X=250880 $Y=91710
X305 3 MASCO__Y24 $T=252495 145110 0 0 $X=252495 $Y=145110
X306 4 MASCO__Y24 $T=266880 91710 0 0 $X=266880 $Y=91710
X307 4 MASCO__Y24 $T=282880 91710 0 0 $X=282880 $Y=91710
X308 4 MASCO__Y24 $T=298880 91710 0 0 $X=298880 $Y=91710
X309 4 MASCO__Y24 $T=314880 91710 0 0 $X=314880 $Y=91710
X310 4 MASCO__Y24 $T=330880 91710 0 0 $X=330880 $Y=91710
.ends MASCO__H1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246551802831                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246551802831 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246551802831

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246551802852                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246551802852 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246551802852

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X4                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X4 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7246551802815 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7246551802815 $T=500 2500 0 0 $X=0 $Y=2000
X2 1 VIATP_C_CDNS_7246551802815 $T=500 4500 0 0 $X=0 $Y=4000
X3 1 VIATP_C_CDNS_7246551802815 $T=500 6500 0 0 $X=0 $Y=6000
X4 1 VIATP_C_CDNS_7246551802815 $T=500 8500 0 0 $X=0 $Y=8000
X5 1 VIATP_C_CDNS_7246551802815 $T=500 10500 0 0 $X=0 $Y=10000
.ends MASCO__X4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X5                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X5 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7246551802815 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7246551802815 $T=500 2500 0 0 $X=0 $Y=2000
X2 1 VIATP_C_CDNS_7246551802815 $T=500 4500 0 0 $X=0 $Y=4000
X3 1 VIATP_C_CDNS_7246551802815 $T=500 6500 0 0 $X=0 $Y=6000
X4 1 VIATP_C_CDNS_7246551802815 $T=500 8500 0 0 $X=0 $Y=8000
X5 1 VIATP_C_CDNS_7246551802815 $T=500 10500 0 0 $X=0 $Y=10000
X6 1 VIATP_C_CDNS_7246551802815 $T=500 12500 0 0 $X=0 $Y=12000
.ends MASCO__X5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X6                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X6 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7246551802815 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7246551802815 $T=500 1500 0 0 $X=0 $Y=1000
X2 1 VIATP_C_CDNS_7246551802815 $T=500 2500 0 0 $X=0 $Y=2000
X3 1 VIATP_C_CDNS_7246551802815 $T=500 3500 0 0 $X=0 $Y=3000
X4 1 VIATP_C_CDNS_7246551802815 $T=500 4500 0 0 $X=0 $Y=4000
X5 1 VIATP_C_CDNS_7246551802815 $T=500 5500 0 0 $X=0 $Y=5000
X6 1 VIATP_C_CDNS_7246551802815 $T=500 6500 0 0 $X=0 $Y=6000
X7 1 VIATP_C_CDNS_7246551802815 $T=500 7500 0 0 $X=0 $Y=7000
X8 1 VIATP_C_CDNS_7246551802815 $T=500 8500 0 0 $X=0 $Y=8000
.ends MASCO__X6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X7                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X7 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7246551802815 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7246551802815 $T=500 1500 0 0 $X=0 $Y=1000
X2 1 VIATP_C_CDNS_7246551802815 $T=500 2500 0 0 $X=0 $Y=2000
X3 1 VIATP_C_CDNS_7246551802815 $T=500 3500 0 0 $X=0 $Y=3000
X4 1 VIATP_C_CDNS_7246551802815 $T=500 4500 0 0 $X=0 $Y=4000
X5 1 VIATP_C_CDNS_7246551802815 $T=500 5500 0 0 $X=0 $Y=5000
X6 1 VIATP_C_CDNS_7246551802815 $T=500 6500 0 0 $X=0 $Y=6000
X7 1 VIATP_C_CDNS_7246551802815 $T=500 7500 0 0 $X=0 $Y=7000
.ends MASCO__X7

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y20                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y20 1
** N=1 EP=1 FDC=0
X0 1 MASCO__X6 $T=0 0 0 0 $X=0 $Y=0
X1 1 MASCO__X6 $T=2000 0 0 0 $X=2000 $Y=0
X2 1 MASCO__X6 $T=4000 0 0 0 $X=4000 $Y=0
X3 1 MASCO__X6 $T=6000 0 0 0 $X=6000 $Y=0
X4 1 MASCO__X6 $T=8000 0 0 0 $X=8000 $Y=0
X5 1 MASCO__X6 $T=10000 0 0 0 $X=10000 $Y=0
X6 1 MASCO__X6 $T=12000 0 0 0 $X=12000 $Y=0
X7 1 MASCO__X6 $T=14000 0 0 0 $X=14000 $Y=0
.ends MASCO__Y20

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y21                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y21 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7246551802831 $T=500 750 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7246551802831 $T=1500 750 0 0 $X=1000 $Y=0
X2 1 VIATP_C_CDNS_7246551802831 $T=2500 750 0 0 $X=2000 $Y=0
X3 1 VIATP_C_CDNS_7246551802831 $T=3500 750 0 0 $X=3000 $Y=0
X4 1 VIATP_C_CDNS_7246551802831 $T=4500 750 0 0 $X=4000 $Y=0
X5 1 VIATP_C_CDNS_7246551802831 $T=5500 750 0 0 $X=5000 $Y=0
X6 1 VIATP_C_CDNS_7246551802831 $T=6500 750 0 0 $X=6000 $Y=0
X7 1 VIATP_C_CDNS_7246551802831 $T=7500 750 0 0 $X=7000 $Y=0
X8 1 VIATP_C_CDNS_7246551802831 $T=8500 750 0 0 $X=8000 $Y=0
X9 1 VIATP_C_CDNS_7246551802831 $T=9500 750 0 0 $X=9000 $Y=0
X10 1 VIATP_C_CDNS_7246551802831 $T=10500 750 0 0 $X=10000 $Y=0
X11 1 VIATP_C_CDNS_7246551802831 $T=11500 750 0 0 $X=11000 $Y=0
.ends MASCO__Y21

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X8                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X8 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7246551802815 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7246551802815 $T=500 2500 0 0 $X=0 $Y=2000
X2 1 VIATP_C_CDNS_7246551802815 $T=500 4500 0 0 $X=0 $Y=4000
X3 1 VIATP_C_CDNS_7246551802815 $T=500 6500 0 0 $X=0 $Y=6000
X4 1 VIATP_C_CDNS_7246551802815 $T=500 8500 0 0 $X=0 $Y=8000
X5 1 VIATP_C_CDNS_7246551802815 $T=500 10500 0 0 $X=0 $Y=10000
X6 1 VIATP_C_CDNS_7246551802815 $T=500 12500 0 0 $X=0 $Y=12000
X7 1 VIATP_C_CDNS_7246551802815 $T=500 14500 0 0 $X=0 $Y=14000
.ends MASCO__X8

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y22                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y22 1
** N=1 EP=1 FDC=0
X0 1 MASCO__X8 $T=0 0 0 0 $X=0 $Y=0
X1 1 MASCO__X8 $T=2000 0 0 0 $X=2000 $Y=0
X2 1 MASCO__X8 $T=4000 0 0 0 $X=4000 $Y=0
X3 1 MASCO__X8 $T=6000 0 0 0 $X=6000 $Y=0
.ends MASCO__Y22

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__P2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__P2 1 2 3 4 5 6
** N=6 EP=6 FDC=370
X0 6 VIATP_C_CDNS_7246551802831 $T=342380 73960 0 0 $X=341880 $Y=73210
X1 6 VIATP_C_CDNS_7246551802831 $T=343380 73960 0 0 $X=342880 $Y=73210
X2 6 VIATP_C_CDNS_7246551802831 $T=344380 73960 0 0 $X=343880 $Y=73210
X3 6 VIATP_C_CDNS_7246551802831 $T=345380 73960 0 0 $X=344880 $Y=73210
X4 6 VIATP_C_CDNS_7246551802831 $T=346380 73960 0 0 $X=345880 $Y=73210
X5 6 VIATP_C_CDNS_7246551802831 $T=372380 73960 0 0 $X=371880 $Y=73210
X6 6 VIATP_C_CDNS_7246551802831 $T=373380 73960 0 0 $X=372880 $Y=73210
X7 6 VIATP_C_CDNS_7246551802831 $T=374380 73960 0 0 $X=373880 $Y=73210
X8 6 VIATP_C_CDNS_7246551802831 $T=375380 73960 0 0 $X=374880 $Y=73210
X9 6 VIATP_C_CDNS_7246551802831 $T=376380 73960 0 0 $X=375880 $Y=73210
X10 6 VIATP_C_CDNS_7246551802831 $T=378380 73960 0 0 $X=377880 $Y=73210
X11 6 VIATP_C_CDNS_7246551802831 $T=379380 73960 0 0 $X=378880 $Y=73210
X12 6 VIATP_C_CDNS_7246551802831 $T=380380 73960 0 0 $X=379880 $Y=73210
X13 6 VIATP_C_CDNS_7246551802831 $T=381380 73960 0 0 $X=380880 $Y=73210
X14 6 VIATP_C_CDNS_7246551802831 $T=382380 73960 0 0 $X=381880 $Y=73210
X15 6 VIATP_C_CDNS_7246551802831 $T=383380 73960 0 0 $X=382880 $Y=73210
X16 6 VIATP_C_CDNS_7246551802831 $T=384380 73960 0 0 $X=383880 $Y=73210
X17 6 VIATP_C_CDNS_7246551802831 $T=385380 73960 0 0 $X=384880 $Y=73210
X18 6 VIATP_C_CDNS_7246551802831 $T=386380 73960 0 0 $X=385880 $Y=73210
X19 6 VIATP_C_CDNS_7246551802831 $T=387380 73960 0 0 $X=386880 $Y=73210
X20 6 VIATP_C_CDNS_7246551802831 $T=388380 73960 0 0 $X=387880 $Y=73210
X21 6 VIATP_C_CDNS_7246551802831 $T=389380 73960 0 0 $X=388880 $Y=73210
X22 6 VIATP_C_CDNS_7246551802831 $T=390380 73960 0 0 $X=389880 $Y=73210
X23 6 VIATP_C_CDNS_7246551802831 $T=391380 73960 0 0 $X=390880 $Y=73210
X24 6 VIATP_C_CDNS_7246551802831 $T=392380 73960 0 0 $X=391880 $Y=73210
X25 6 VIATP_C_CDNS_7246551802831 $T=393380 73960 0 0 $X=392880 $Y=73210
X26 6 VIATP_C_CDNS_7246551802831 $T=394380 73960 0 0 $X=393880 $Y=73210
X27 6 VIATP_C_CDNS_7246551802831 $T=395380 73960 0 0 $X=394880 $Y=73210
X28 6 VIATP_C_CDNS_7246551802831 $T=396380 73960 0 0 $X=395880 $Y=73210
X29 6 VIATP_C_CDNS_7246551802831 $T=397380 73960 0 0 $X=396880 $Y=73210
X30 6 VIATP_C_CDNS_7246551802831 $T=398380 73960 0 0 $X=397880 $Y=73210
X31 6 VIATP_C_CDNS_7246551802831 $T=399380 73960 0 0 $X=398880 $Y=73210
X32 6 VIATP_C_CDNS_7246551802831 $T=400380 73960 0 0 $X=399880 $Y=73210
X33 6 VIATP_C_CDNS_7246551802831 $T=401380 73960 0 0 $X=400880 $Y=73210
X34 6 VIATP_C_CDNS_7246551802831 $T=402380 73960 0 0 $X=401880 $Y=73210
X35 6 VIATP_C_CDNS_7246551802833 $T=386380 102330 0 0 $X=385880 $Y=101710
X36 6 VIATP_C_CDNS_7246551802833 $T=387380 102330 0 0 $X=386880 $Y=101710
X37 6 VIATP_C_CDNS_7246551802833 $T=388380 102330 0 0 $X=387880 $Y=101710
X38 6 VIATP_C_CDNS_7246551802833 $T=389380 102330 0 0 $X=388880 $Y=101710
X39 6 VIATP_C_CDNS_7246551802833 $T=390380 102330 0 0 $X=389880 $Y=101710
X40 6 VIATP_C_CDNS_7246551802833 $T=391380 102330 0 0 $X=390880 $Y=101710
X41 6 VIATP_C_CDNS_7246551802833 $T=392380 102330 0 0 $X=391880 $Y=101710
X42 6 VIATP_C_CDNS_7246551802833 $T=393380 102330 0 0 $X=392880 $Y=101710
X43 6 VIATP_C_CDNS_7246551802833 $T=394380 102330 0 0 $X=393880 $Y=101710
X44 6 VIATP_C_CDNS_7246551802833 $T=395380 102330 0 0 $X=394880 $Y=101710
X45 6 VIATP_C_CDNS_7246551802833 $T=396380 102330 0 0 $X=395880 $Y=101710
X46 6 VIATP_C_CDNS_7246551802833 $T=397380 102330 0 0 $X=396880 $Y=101710
X47 6 VIATP_C_CDNS_7246551802833 $T=398380 102330 0 0 $X=397880 $Y=101710
X48 6 VIATP_C_CDNS_7246551802833 $T=399380 102330 0 0 $X=398880 $Y=101710
X49 6 VIATP_C_CDNS_7246551802833 $T=400380 102330 0 0 $X=399880 $Y=101710
X50 6 VIATP_C_CDNS_7246551802833 $T=401380 102330 0 0 $X=400880 $Y=101710
X51 6 VIATP_C_CDNS_7246551802833 $T=402380 102330 0 0 $X=401880 $Y=101710
X52 6 VIATP_C_CDNS_7246551802850 $T=403810 102330 0 0 $X=402880 $Y=101710
X53 6 VIATP_C_CDNS_7246551802851 $T=232950 75210 0 0 $X=232020 $Y=74710
X54 6 VIATP_C_CDNS_7246551802851 $T=232950 76210 0 0 $X=232020 $Y=75710
X55 6 VIATP_C_CDNS_7246551802851 $T=232950 77210 0 0 $X=232020 $Y=76710
X56 6 VIATP_C_CDNS_7246551802851 $T=232950 78210 0 0 $X=232020 $Y=77710
X57 6 VIATP_C_CDNS_7246551802851 $T=232950 79210 0 0 $X=232020 $Y=78710
X58 6 VIATP_C_CDNS_7246551802851 $T=232950 80210 0 0 $X=232020 $Y=79710
X59 6 VIATP_C_CDNS_7246551802851 $T=232950 81210 0 0 $X=232020 $Y=80710
X60 6 VIATP_C_CDNS_7246551802851 $T=232950 82210 0 0 $X=232020 $Y=81710
X61 6 VIATP_C_CDNS_7246551802851 $T=232950 83210 0 0 $X=232020 $Y=82710
X62 6 VIATP_C_CDNS_7246551802851 $T=232950 84210 0 0 $X=232020 $Y=83710
X63 6 VIATP_C_CDNS_7246551802851 $T=232950 85210 0 0 $X=232020 $Y=84710
X64 6 VIATP_C_CDNS_7246551802851 $T=232950 86210 0 0 $X=232020 $Y=85710
X65 6 VIATP_C_CDNS_7246551802851 $T=232950 87210 0 0 $X=232020 $Y=86710
X66 6 VIATP_C_CDNS_7246551802851 $T=232950 88210 0 0 $X=232020 $Y=87710
X67 6 VIATP_C_CDNS_7246551802851 $T=232950 89210 0 0 $X=232020 $Y=88710
X68 6 VIATP_C_CDNS_7246551802851 $T=232950 90210 0 0 $X=232020 $Y=89710
X69 6 VIATP_C_CDNS_7246551802851 $T=232950 91210 0 0 $X=232020 $Y=90710
X70 6 VIATP_C_CDNS_7246551802851 $T=403810 75210 0 0 $X=402880 $Y=74710
X71 6 VIATP_C_CDNS_7246551802851 $T=403810 76210 0 0 $X=402880 $Y=75710
X72 6 VIATP_C_CDNS_7246551802851 $T=403810 77210 0 0 $X=402880 $Y=76710
X73 6 VIATP_C_CDNS_7246551802851 $T=403810 78210 0 0 $X=402880 $Y=77710
X74 6 VIATP_C_CDNS_7246551802851 $T=403810 79210 0 0 $X=402880 $Y=78710
X75 6 VIATP_C_CDNS_7246551802851 $T=403810 80210 0 0 $X=402880 $Y=79710
X76 6 VIATP_C_CDNS_7246551802851 $T=403810 81210 0 0 $X=402880 $Y=80710
X77 6 VIATP_C_CDNS_7246551802851 $T=403810 82210 0 0 $X=402880 $Y=81710
X78 6 VIATP_C_CDNS_7246551802851 $T=403810 83210 0 0 $X=402880 $Y=82710
X79 6 VIATP_C_CDNS_7246551802851 $T=403810 84210 0 0 $X=402880 $Y=83710
X80 6 VIATP_C_CDNS_7246551802851 $T=403810 85210 0 0 $X=402880 $Y=84710
X81 6 VIATP_C_CDNS_7246551802851 $T=403810 86210 0 0 $X=402880 $Y=85710
X82 6 VIATP_C_CDNS_7246551802851 $T=403810 87210 0 0 $X=402880 $Y=86710
X83 6 VIATP_C_CDNS_7246551802851 $T=403810 88210 0 0 $X=402880 $Y=87710
X84 6 VIATP_C_CDNS_7246551802851 $T=403810 89210 0 0 $X=402880 $Y=88710
X85 6 VIATP_C_CDNS_7246551802851 $T=403810 90210 0 0 $X=402880 $Y=89710
X86 6 VIATP_C_CDNS_7246551802851 $T=403810 91210 0 0 $X=402880 $Y=90710
X87 6 VIATP_C_CDNS_7246551802851 $T=403810 92210 0 0 $X=402880 $Y=91710
X88 6 VIATP_C_CDNS_7246551802851 $T=403810 93210 0 0 $X=402880 $Y=92710
X89 6 VIATP_C_CDNS_7246551802851 $T=403810 94210 0 0 $X=402880 $Y=93710
X90 6 VIATP_C_CDNS_7246551802851 $T=403810 95210 0 0 $X=402880 $Y=94710
X91 6 VIATP_C_CDNS_7246551802851 $T=403810 96210 0 0 $X=402880 $Y=95710
X92 6 VIATP_C_CDNS_7246551802851 $T=403810 97210 0 0 $X=402880 $Y=96710
X93 6 VIATP_C_CDNS_7246551802851 $T=403810 98210 0 0 $X=402880 $Y=97710
X94 6 VIATP_C_CDNS_7246551802851 $T=403810 99210 0 0 $X=402880 $Y=98710
X95 6 VIATP_C_CDNS_7246551802851 $T=403810 100210 0 0 $X=402880 $Y=99710
X96 6 VIATP_C_CDNS_7246551802851 $T=403810 101210 0 0 $X=402880 $Y=100710
X97 6 VIATP_C_CDNS_7246551802852 $T=232950 73960 0 0 $X=232020 $Y=73210
X98 6 VIATP_C_CDNS_7246551802852 $T=403810 73960 0 0 $X=402880 $Y=73210
X99 6 VIATP_C_CDNS_7246551802854 $T=377440 75210 0 0 $X=377000 $Y=74710
X100 6 VIATP_C_CDNS_7246551802854 $T=377440 76210 0 0 $X=377000 $Y=75710
X101 6 VIATP_C_CDNS_7246551802854 $T=377440 77210 0 0 $X=377000 $Y=76710
X102 6 VIATP_C_CDNS_7246551802854 $T=377440 78210 0 0 $X=377000 $Y=77710
X103 6 VIATP_C_CDNS_7246551802854 $T=377440 79210 0 0 $X=377000 $Y=78710
X104 6 VIATP_C_CDNS_7246551802854 $T=377440 80210 0 0 $X=377000 $Y=79710
X105 6 VIATP_C_CDNS_7246551802854 $T=377440 81210 0 0 $X=377000 $Y=80710
X106 6 VIATP_C_CDNS_7246551802854 $T=377440 82210 0 0 $X=377000 $Y=81710
X107 6 VIATP_C_CDNS_7246551802854 $T=377440 83210 0 0 $X=377000 $Y=82710
X108 6 VIATP_C_CDNS_7246551802854 $T=377440 84210 0 0 $X=377000 $Y=83710
X109 6 VIATP_C_CDNS_7246551802854 $T=377440 85210 0 0 $X=377000 $Y=84710
X110 6 VIATP_C_CDNS_7246551802854 $T=377440 86210 0 0 $X=377000 $Y=85710
X111 6 VIATP_C_CDNS_7246551802854 $T=377440 87210 0 0 $X=377000 $Y=86710
X112 6 VIATP_C_CDNS_7246551802854 $T=377440 88210 0 0 $X=377000 $Y=87710
X113 6 VIATP_C_CDNS_7246551802854 $T=377440 89210 0 0 $X=377000 $Y=88710
X114 6 VIATP_C_CDNS_7246551802854 $T=377440 90210 0 0 $X=377000 $Y=89710
X115 6 VIATP_C_CDNS_7246551802854 $T=377440 91210 0 0 $X=377000 $Y=90710
X116 6 MASCO__X4 $T=385880 89710 0 0 $X=385880 $Y=89710
X117 6 MASCO__X4 $T=387880 89710 0 0 $X=387880 $Y=89710
X118 6 MASCO__X4 $T=389880 89710 0 0 $X=389880 $Y=89710
X119 6 MASCO__X4 $T=391880 89710 0 0 $X=391880 $Y=89710
X120 6 MASCO__X4 $T=393880 89710 0 0 $X=393880 $Y=89710
X121 6 MASCO__X4 $T=395880 89710 0 0 $X=395880 $Y=89710
X122 6 MASCO__X4 $T=397880 89710 0 0 $X=397880 $Y=89710
X123 6 MASCO__X4 $T=399880 89710 0 0 $X=399880 $Y=89710
X124 6 MASCO__X4 $T=401880 89710 0 0 $X=401880 $Y=89710
X125 6 MASCO__X5 $T=385880 75710 0 0 $X=385880 $Y=75710
X126 6 MASCO__X5 $T=387880 75710 0 0 $X=387880 $Y=75710
X127 6 MASCO__X5 $T=389880 75710 0 0 $X=389880 $Y=75710
X128 6 MASCO__X5 $T=391880 75710 0 0 $X=391880 $Y=75710
X129 6 MASCO__X5 $T=393880 75710 0 0 $X=393880 $Y=75710
X130 6 MASCO__X5 $T=395880 75710 0 0 $X=395880 $Y=75710
X131 6 MASCO__X5 $T=397880 75710 0 0 $X=397880 $Y=75710
X132 6 MASCO__X5 $T=399880 75710 0 0 $X=399880 $Y=75710
X133 6 MASCO__X5 $T=401880 75710 0 0 $X=401880 $Y=75710
X134 6 MASCO__X6 $T=348880 74710 0 0 $X=348880 $Y=74710
X135 6 MASCO__X6 $T=350880 74710 0 0 $X=350880 $Y=74710
X136 6 MASCO__X6 $T=352880 74710 0 0 $X=352880 $Y=74710
X137 6 MASCO__X6 $T=354880 74710 0 0 $X=354880 $Y=74710
X138 6 MASCO__X6 $T=356880 74710 0 0 $X=356880 $Y=74710
X139 6 MASCO__X6 $T=358880 74710 0 0 $X=358880 $Y=74710
X140 6 MASCO__X6 $T=360880 74710 0 0 $X=360880 $Y=74710
X141 6 MASCO__X6 $T=362880 74710 0 0 $X=362880 $Y=74710
X142 6 MASCO__X6 $T=364880 74710 0 0 $X=364880 $Y=74710
X143 6 MASCO__X6 $T=366880 74710 0 0 $X=366880 $Y=74710
X144 6 MASCO__X6 $T=368880 74710 0 0 $X=368880 $Y=74710
X145 6 MASCO__X6 $T=370880 74710 0 0 $X=370880 $Y=74710
X146 6 MASCO__X6 $T=372880 74710 0 0 $X=372880 $Y=74710
X147 6 MASCO__X6 $T=374880 74710 0 0 $X=374880 $Y=74710
X148 6 MASCO__X6 $T=378880 74710 0 0 $X=378880 $Y=74710
X149 6 MASCO__X6 $T=380880 74710 0 0 $X=380880 $Y=74710
X150 6 MASCO__X6 $T=382880 74710 0 0 $X=382880 $Y=74710
X151 6 MASCO__X6 $T=384880 74710 0 0 $X=384880 $Y=74710
X152 6 MASCO__X6 $T=386880 74710 0 0 $X=386880 $Y=74710
X153 6 MASCO__X6 $T=388880 74710 0 0 $X=388880 $Y=74710
X154 6 MASCO__X6 $T=390880 74710 0 0 $X=390880 $Y=74710
X155 6 MASCO__X6 $T=392880 74710 0 0 $X=392880 $Y=74710
X156 6 MASCO__X6 $T=394880 74710 0 0 $X=394880 $Y=74710
X157 6 MASCO__X6 $T=396880 74710 0 0 $X=396880 $Y=74710
X158 6 MASCO__X6 $T=398880 74710 0 0 $X=398880 $Y=74710
X159 6 MASCO__X6 $T=400880 74710 0 0 $X=400880 $Y=74710
X160 6 MASCO__X7 $T=234880 83710 0 0 $X=234880 $Y=83710
X161 6 MASCO__X7 $T=236880 83710 0 0 $X=236880 $Y=83710
X162 6 MASCO__X7 $T=238880 83710 0 0 $X=238880 $Y=83710
X163 6 MASCO__X7 $T=240880 83710 0 0 $X=240880 $Y=83710
X164 6 MASCO__X7 $T=242880 83710 0 0 $X=242880 $Y=83710
X165 6 MASCO__X7 $T=244880 83710 0 0 $X=244880 $Y=83710
X166 6 MASCO__X7 $T=246880 83710 0 0 $X=246880 $Y=83710
X167 6 MASCO__X7 $T=248880 83710 0 0 $X=248880 $Y=83710
X168 6 MASCO__X7 $T=250880 83710 0 0 $X=250880 $Y=83710
X169 6 MASCO__X7 $T=252880 83710 0 0 $X=252880 $Y=83710
X170 6 MASCO__X7 $T=254880 83710 0 0 $X=254880 $Y=83710
X171 6 MASCO__X7 $T=256880 83710 0 0 $X=256880 $Y=83710
X172 6 MASCO__X7 $T=258880 83710 0 0 $X=258880 $Y=83710
X173 6 MASCO__X7 $T=260880 83710 0 0 $X=260880 $Y=83710
X174 6 MASCO__X7 $T=262880 83710 0 0 $X=262880 $Y=83710
X175 6 MASCO__X7 $T=264880 83710 0 0 $X=264880 $Y=83710
X176 6 MASCO__X7 $T=266880 83710 0 0 $X=266880 $Y=83710
X177 6 MASCO__X7 $T=268880 83710 0 0 $X=268880 $Y=83710
X178 6 MASCO__X7 $T=270880 83710 0 0 $X=270880 $Y=83710
X179 6 MASCO__X7 $T=272880 83710 0 0 $X=272880 $Y=83710
X180 6 MASCO__X7 $T=274880 83710 0 0 $X=274880 $Y=83710
X181 6 MASCO__X7 $T=276880 83710 0 0 $X=276880 $Y=83710
X182 6 MASCO__X7 $T=278880 83710 0 0 $X=278880 $Y=83710
X183 6 MASCO__X7 $T=280880 83710 0 0 $X=280880 $Y=83710
X184 6 MASCO__X7 $T=282880 83710 0 0 $X=282880 $Y=83710
X185 6 MASCO__X7 $T=284880 83710 0 0 $X=284880 $Y=83710
X186 6 MASCO__X7 $T=286880 83710 0 0 $X=286880 $Y=83710
X187 6 MASCO__X7 $T=288880 83710 0 0 $X=288880 $Y=83710
X188 6 MASCO__X7 $T=290880 83710 0 0 $X=290880 $Y=83710
X189 6 MASCO__X7 $T=292880 83710 0 0 $X=292880 $Y=83710
X190 6 MASCO__X7 $T=294880 83710 0 0 $X=294880 $Y=83710
X191 6 MASCO__X7 $T=296880 83710 0 0 $X=296880 $Y=83710
X192 6 MASCO__X7 $T=298880 83710 0 0 $X=298880 $Y=83710
X193 6 MASCO__X7 $T=300880 83710 0 0 $X=300880 $Y=83710
X194 6 MASCO__X7 $T=302880 83710 0 0 $X=302880 $Y=83710
X195 6 MASCO__X7 $T=304880 83710 0 0 $X=304880 $Y=83710
X196 6 MASCO__X7 $T=306880 83710 0 0 $X=306880 $Y=83710
X197 6 MASCO__X7 $T=308880 83710 0 0 $X=308880 $Y=83710
X198 6 MASCO__X7 $T=310880 83710 0 0 $X=310880 $Y=83710
X199 6 MASCO__X7 $T=312880 83710 0 0 $X=312880 $Y=83710
X200 6 MASCO__X7 $T=314880 83710 0 0 $X=314880 $Y=83710
X201 6 MASCO__X7 $T=316880 83710 0 0 $X=316880 $Y=83710
X202 6 MASCO__X7 $T=318880 83710 0 0 $X=318880 $Y=83710
X203 6 MASCO__X7 $T=320880 83710 0 0 $X=320880 $Y=83710
X204 6 MASCO__X7 $T=322880 83710 0 0 $X=322880 $Y=83710
X205 6 MASCO__X7 $T=324880 83710 0 0 $X=324880 $Y=83710
X206 6 MASCO__X7 $T=326880 83710 0 0 $X=326880 $Y=83710
X207 6 MASCO__X7 $T=328880 83710 0 0 $X=328880 $Y=83710
X208 6 MASCO__X7 $T=330880 83710 0 0 $X=330880 $Y=83710
X209 6 MASCO__X7 $T=332880 83710 0 0 $X=332880 $Y=83710
X210 6 MASCO__X7 $T=334880 83710 0 0 $X=334880 $Y=83710
X211 6 MASCO__X7 $T=336880 83710 0 0 $X=336880 $Y=83710
X212 6 MASCO__X7 $T=338880 83710 0 0 $X=338880 $Y=83710
X213 6 MASCO__X7 $T=340880 83710 0 0 $X=340880 $Y=83710
X214 6 MASCO__X7 $T=342880 83710 0 0 $X=342880 $Y=83710
X215 6 MASCO__X7 $T=344880 83710 0 0 $X=344880 $Y=83710
X216 6 MASCO__X7 $T=348880 83710 0 0 $X=348880 $Y=83710
X217 6 MASCO__X7 $T=350880 83710 0 0 $X=350880 $Y=83710
X218 6 MASCO__X7 $T=352880 83710 0 0 $X=352880 $Y=83710
X219 6 MASCO__X7 $T=354880 83710 0 0 $X=354880 $Y=83710
X220 6 MASCO__X7 $T=356880 83710 0 0 $X=356880 $Y=83710
X221 6 MASCO__X7 $T=358880 83710 0 0 $X=358880 $Y=83710
X222 6 MASCO__X7 $T=360880 83710 0 0 $X=360880 $Y=83710
X223 6 MASCO__X7 $T=362880 83710 0 0 $X=362880 $Y=83710
X224 6 MASCO__X7 $T=364880 83710 0 0 $X=364880 $Y=83710
X225 6 MASCO__X7 $T=366880 83710 0 0 $X=366880 $Y=83710
X226 6 MASCO__X7 $T=368880 83710 0 0 $X=368880 $Y=83710
X227 6 MASCO__X7 $T=370880 83710 0 0 $X=370880 $Y=83710
X228 6 MASCO__X7 $T=372880 83710 0 0 $X=372880 $Y=83710
X229 6 MASCO__X7 $T=374880 83710 0 0 $X=374880 $Y=83710
X230 6 MASCO__X7 $T=378880 83710 0 0 $X=378880 $Y=83710
X231 6 MASCO__X7 $T=380880 83710 0 0 $X=380880 $Y=83710
X232 6 MASCO__X7 $T=382880 83710 0 0 $X=382880 $Y=83710
X233 6 MASCO__X7 $T=384880 83710 0 0 $X=384880 $Y=83710
X234 6 MASCO__Y20 $T=234880 74710 0 0 $X=234880 $Y=74710
X235 6 MASCO__Y20 $T=250880 74710 0 0 $X=250880 $Y=74710
X236 6 MASCO__Y20 $T=266880 74710 0 0 $X=266880 $Y=74710
X237 6 MASCO__Y20 $T=282880 74710 0 0 $X=282880 $Y=74710
X238 6 MASCO__Y20 $T=298880 74710 0 0 $X=298880 $Y=74710
X239 6 MASCO__Y20 $T=314880 74710 0 0 $X=314880 $Y=74710
X240 6 MASCO__Y20 $T=330880 74710 0 0 $X=330880 $Y=74710
X241 6 MASCO__Y20 $T=386880 83710 0 0 $X=386880 $Y=83710
X242 6 MASCO__Y20 $T=386880 92710 0 0 $X=386880 $Y=92710
X243 6 MASCO__Y21 $T=233880 73210 0 0 $X=233880 $Y=73210
X244 6 MASCO__Y21 $T=245880 73210 0 0 $X=245880 $Y=73210
X245 6 MASCO__Y21 $T=257880 73210 0 0 $X=257880 $Y=73210
X246 6 MASCO__Y21 $T=269880 73210 0 0 $X=269880 $Y=73210
X247 6 MASCO__Y21 $T=281880 73210 0 0 $X=281880 $Y=73210
X248 6 MASCO__Y21 $T=293880 73210 0 0 $X=293880 $Y=73210
X249 6 MASCO__Y21 $T=305880 73210 0 0 $X=305880 $Y=73210
X250 6 MASCO__Y21 $T=317880 73210 0 0 $X=317880 $Y=73210
X251 6 MASCO__Y21 $T=329880 73210 0 0 $X=329880 $Y=73210
X252 6 MASCO__Y21 $T=347880 73210 0 0 $X=347880 $Y=73210
X253 6 MASCO__Y21 $T=359880 73210 0 0 $X=359880 $Y=73210
X254 6 MASCO__Y22 $T=233880 75710 0 0 $X=233880 $Y=75710
X255 6 MASCO__Y22 $T=241880 75710 0 0 $X=241880 $Y=75710
X256 6 MASCO__Y22 $T=249880 75710 0 0 $X=249880 $Y=75710
X257 6 MASCO__Y22 $T=257880 75710 0 0 $X=257880 $Y=75710
X258 6 MASCO__Y22 $T=265880 75710 0 0 $X=265880 $Y=75710
X259 6 MASCO__Y22 $T=273880 75710 0 0 $X=273880 $Y=75710
X260 6 MASCO__Y22 $T=281880 75710 0 0 $X=281880 $Y=75710
X261 6 MASCO__Y22 $T=289880 75710 0 0 $X=289880 $Y=75710
X262 6 MASCO__Y22 $T=297880 75710 0 0 $X=297880 $Y=75710
X263 6 MASCO__Y22 $T=305880 75710 0 0 $X=305880 $Y=75710
X264 6 MASCO__Y22 $T=313880 75710 0 0 $X=313880 $Y=75710
X265 6 MASCO__Y22 $T=321880 75710 0 0 $X=321880 $Y=75710
X266 6 MASCO__Y22 $T=329880 75710 0 0 $X=329880 $Y=75710
X267 6 MASCO__Y22 $T=337880 75710 0 0 $X=337880 $Y=75710
X268 6 MASCO__Y22 $T=345880 75710 0 0 $X=345880 $Y=75710
X269 6 MASCO__Y22 $T=353880 75710 0 0 $X=353880 $Y=75710
X270 6 MASCO__Y22 $T=361880 75710 0 0 $X=361880 $Y=75710
X271 6 MASCO__Y22 $T=369880 75710 0 0 $X=369880 $Y=75710
X272 6 MASCO__Y22 $T=377880 75710 0 0 $X=377880 $Y=75710
C0 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=11155 $Y=41445 $dt=11
C1 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=11155 $Y=47485 $dt=11
C2 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=11155 $Y=53525 $dt=11
C3 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=11155 $Y=59565 $dt=11
C4 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=11155 $Y=65605 $dt=11
C5 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=11155 $Y=71645 $dt=11
C6 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=11155 $Y=77685 $dt=11
C7 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=11155 $Y=83725 $dt=11
C8 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=11155 $Y=89765 $dt=11
C9 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=11155 $Y=95805 $dt=11
C10 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=12135 $Y=10115 $dt=11
C11 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=12135 $Y=21815 $dt=11
C12 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=18175 $Y=10115 $dt=11
C13 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=18175 $Y=21815 $dt=11
C14 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=22855 $Y=41445 $dt=11
C15 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=22855 $Y=47485 $dt=11
C16 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=22855 $Y=53525 $dt=11
C17 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=22855 $Y=59565 $dt=11
C18 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=22855 $Y=65605 $dt=11
C19 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=22855 $Y=71645 $dt=11
C20 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=22855 $Y=77685 $dt=11
C21 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=22855 $Y=83725 $dt=11
C22 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=22855 $Y=89765 $dt=11
C23 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=22855 $Y=95805 $dt=11
C24 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=24215 $Y=10115 $dt=11
C25 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=24215 $Y=21815 $dt=11
C26 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=30255 $Y=10115 $dt=11
C27 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=30255 $Y=21815 $dt=11
C28 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=34555 $Y=41445 $dt=11
C29 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=34555 $Y=47485 $dt=11
C30 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=34555 $Y=53525 $dt=11
C31 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=34555 $Y=59565 $dt=11
C32 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=34555 $Y=65605 $dt=11
C33 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=34555 $Y=71645 $dt=11
C34 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=34555 $Y=77685 $dt=11
C35 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=34555 $Y=83725 $dt=11
C36 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=34555 $Y=89765 $dt=11
C37 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=34555 $Y=95805 $dt=11
C38 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=36295 $Y=10115 $dt=11
C39 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=36295 $Y=21815 $dt=11
C40 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=42335 $Y=10115 $dt=11
C41 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=42335 $Y=21815 $dt=11
C42 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=46255 $Y=41445 $dt=11
C43 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=46255 $Y=47485 $dt=11
C44 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=46255 $Y=53525 $dt=11
C45 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=46255 $Y=59565 $dt=11
C46 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=46255 $Y=65605 $dt=11
C47 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=46255 $Y=71645 $dt=11
C48 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=46255 $Y=77685 $dt=11
C49 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=46255 $Y=83725 $dt=11
C50 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=46255 $Y=89765 $dt=11
C51 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=46255 $Y=95805 $dt=11
C52 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=48375 $Y=10115 $dt=11
C53 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=48375 $Y=21815 $dt=11
C54 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=54415 $Y=10115 $dt=11
C55 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=54415 $Y=21815 $dt=11
C56 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=57955 $Y=41445 $dt=11
C57 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=57955 $Y=47485 $dt=11
C58 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=57955 $Y=53525 $dt=11
C59 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=57955 $Y=59565 $dt=11
C60 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=57955 $Y=65605 $dt=11
C61 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=57955 $Y=71645 $dt=11
C62 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=57955 $Y=77685 $dt=11
C63 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=57955 $Y=83725 $dt=11
C64 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=57955 $Y=89765 $dt=11
C65 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=57955 $Y=95805 $dt=11
C66 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=60455 $Y=10115 $dt=11
C67 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=60455 $Y=21815 $dt=11
C68 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=66495 $Y=10115 $dt=11
C69 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=66495 $Y=21815 $dt=11
C70 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=69655 $Y=41445 $dt=11
C71 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=69655 $Y=47485 $dt=11
C72 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=69655 $Y=53525 $dt=11
C73 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=69655 $Y=59565 $dt=11
C74 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=69655 $Y=65605 $dt=11
C75 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=69655 $Y=71645 $dt=11
C76 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=69655 $Y=77685 $dt=11
C77 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=69655 $Y=83725 $dt=11
C78 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=69655 $Y=89765 $dt=11
C79 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=69655 $Y=95805 $dt=11
C80 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=72535 $Y=10115 $dt=11
C81 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=72535 $Y=21815 $dt=11
C82 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=78575 $Y=10115 $dt=11
C83 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=78575 $Y=21815 $dt=11
C84 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=81355 $Y=41445 $dt=11
C85 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=81355 $Y=47485 $dt=11
C86 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=81355 $Y=53525 $dt=11
C87 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=81355 $Y=59565 $dt=11
C88 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=81355 $Y=65605 $dt=11
C89 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=81355 $Y=71645 $dt=11
C90 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=81355 $Y=77685 $dt=11
C91 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=81355 $Y=83725 $dt=11
C92 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=81355 $Y=89765 $dt=11
C93 2 5 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=81355 $Y=95805 $dt=11
C94 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=84615 $Y=10115 $dt=11
C95 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=84615 $Y=21815 $dt=11
C96 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=90655 $Y=10115 $dt=11
C97 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=90655 $Y=21815 $dt=11
C98 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=96695 $Y=10115 $dt=11
C99 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=96695 $Y=21815 $dt=11
C100 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=96990 $Y=37085 $dt=11
C101 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=96990 $Y=48785 $dt=11
C102 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=96990 $Y=60485 $dt=11
C103 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=102735 $Y=10115 $dt=11
C104 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=102735 $Y=21815 $dt=11
C105 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=103030 $Y=37085 $dt=11
C106 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=103030 $Y=48785 $dt=11
C107 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=103030 $Y=60485 $dt=11
C108 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=108775 $Y=10115 $dt=11
C109 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=108775 $Y=21815 $dt=11
C110 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=109070 $Y=37085 $dt=11
C111 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=109070 $Y=48785 $dt=11
C112 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=109070 $Y=60485 $dt=11
C113 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=114815 $Y=10115 $dt=11
C114 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=114815 $Y=21815 $dt=11
C115 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=115110 $Y=37085 $dt=11
C116 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=115110 $Y=48785 $dt=11
C117 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=115110 $Y=60485 $dt=11
C118 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=118085 $Y=79030 $dt=11
C119 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=118085 $Y=90730 $dt=11
C120 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=120855 $Y=10115 $dt=11
C121 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=120855 $Y=21815 $dt=11
C122 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=121150 $Y=37085 $dt=11
C123 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=121150 $Y=48785 $dt=11
C124 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=121150 $Y=60485 $dt=11
C125 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=124125 $Y=79030 $dt=11
C126 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=124125 $Y=90730 $dt=11
C127 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=126895 $Y=10115 $dt=11
C128 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=126895 $Y=21815 $dt=11
C129 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=127190 $Y=37085 $dt=11
C130 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=127190 $Y=48785 $dt=11
C131 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=127190 $Y=60485 $dt=11
C132 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=130165 $Y=79030 $dt=11
C133 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=130165 $Y=90730 $dt=11
C134 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=132935 $Y=10115 $dt=11
C135 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=132935 $Y=21815 $dt=11
C136 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=133230 $Y=37085 $dt=11
C137 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=133230 $Y=48785 $dt=11
C138 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=133230 $Y=60485 $dt=11
C139 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=136205 $Y=79030 $dt=11
C140 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=136205 $Y=90730 $dt=11
C141 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=138975 $Y=10115 $dt=11
C142 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=138975 $Y=21815 $dt=11
C143 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=139270 $Y=37085 $dt=11
C144 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=139270 $Y=48785 $dt=11
C145 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=139270 $Y=60485 $dt=11
C146 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=142245 $Y=79030 $dt=11
C147 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=142245 $Y=90730 $dt=11
C148 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=145015 $Y=10115 $dt=11
C149 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=145015 $Y=21815 $dt=11
C150 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=145310 $Y=37085 $dt=11
C151 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=145310 $Y=48785 $dt=11
C152 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=145310 $Y=60485 $dt=11
C153 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=148285 $Y=79030 $dt=11
C154 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=148285 $Y=90730 $dt=11
C155 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=151055 $Y=10115 $dt=11
C156 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=151055 $Y=21815 $dt=11
C157 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=151350 $Y=37085 $dt=11
C158 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=151350 $Y=48785 $dt=11
C159 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=151350 $Y=60485 $dt=11
C160 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=154325 $Y=79030 $dt=11
C161 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=154325 $Y=90730 $dt=11
C162 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=157095 $Y=10115 $dt=11
C163 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=157095 $Y=21815 $dt=11
C164 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=157390 $Y=37085 $dt=11
C165 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=157390 $Y=48785 $dt=11
C166 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=157390 $Y=60485 $dt=11
C167 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=160365 $Y=79030 $dt=11
C168 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=160365 $Y=90730 $dt=11
C169 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=163135 $Y=10115 $dt=11
C170 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=163135 $Y=21815 $dt=11
C171 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=163430 $Y=37085 $dt=11
C172 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=163430 $Y=48785 $dt=11
C173 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=163430 $Y=60485 $dt=11
C174 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=166405 $Y=79030 $dt=11
C175 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=166405 $Y=90730 $dt=11
C176 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=169175 $Y=10115 $dt=11
C177 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=169175 $Y=21815 $dt=11
C178 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=169470 $Y=37085 $dt=11
C179 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=169470 $Y=48785 $dt=11
C180 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=169470 $Y=60485 $dt=11
C181 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=172445 $Y=79030 $dt=11
C182 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=172445 $Y=90730 $dt=11
C183 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=175215 $Y=10115 $dt=11
C184 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=175215 $Y=21815 $dt=11
C185 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=175510 $Y=37085 $dt=11
C186 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=175510 $Y=48785 $dt=11
C187 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=175510 $Y=60485 $dt=11
C188 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=178485 $Y=79030 $dt=11
C189 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=178485 $Y=90730 $dt=11
C190 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=181255 $Y=10115 $dt=11
C191 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=181255 $Y=21815 $dt=11
C192 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=181550 $Y=37085 $dt=11
C193 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=181550 $Y=48785 $dt=11
C194 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=181550 $Y=60485 $dt=11
C195 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=187295 $Y=10115 $dt=11
C196 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=187295 $Y=21815 $dt=11
C197 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=187590 $Y=37085 $dt=11
C198 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=187590 $Y=48785 $dt=11
C199 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=187590 $Y=60485 $dt=11
C200 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=193335 $Y=10115 $dt=11
C201 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=193335 $Y=21815 $dt=11
C202 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=193630 $Y=37085 $dt=11
C203 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=193630 $Y=48785 $dt=11
C204 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=193630 $Y=60485 $dt=11
C205 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=199375 $Y=10115 $dt=11
C206 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=199375 $Y=21815 $dt=11
C207 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=199670 $Y=37085 $dt=11
C208 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=199670 $Y=48785 $dt=11
C209 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=199670 $Y=60485 $dt=11
C210 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=205415 $Y=10115 $dt=11
C211 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=205415 $Y=21815 $dt=11
C212 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=205710 $Y=37085 $dt=11
C213 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=205710 $Y=48785 $dt=11
C214 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=205710 $Y=60485 $dt=11
C215 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=211455 $Y=10115 $dt=11
C216 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=211455 $Y=21815 $dt=11
C217 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=211750 $Y=37085 $dt=11
C218 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=211750 $Y=48785 $dt=11
C219 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=211750 $Y=60485 $dt=11
C220 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=217495 $Y=10115 $dt=11
C221 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=217495 $Y=21815 $dt=11
C222 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=217790 $Y=37085 $dt=11
C223 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=217790 $Y=48785 $dt=11
C224 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=217790 $Y=60485 $dt=11
C225 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=223535 $Y=10115 $dt=11
C226 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=223535 $Y=21815 $dt=11
C227 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=223830 $Y=37085 $dt=11
C228 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=223830 $Y=48785 $dt=11
C229 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=223830 $Y=60485 $dt=11
C230 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=229575 $Y=10115 $dt=11
C231 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=229575 $Y=21815 $dt=11
C232 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=229870 $Y=37085 $dt=11
C233 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=229870 $Y=48785 $dt=11
C234 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=229870 $Y=60485 $dt=11
C235 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=235615 $Y=10115 $dt=11
C236 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=235615 $Y=21815 $dt=11
C237 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=235910 $Y=37085 $dt=11
C238 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=235910 $Y=48785 $dt=11
C239 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=235910 $Y=60485 $dt=11
C240 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=241655 $Y=10115 $dt=11
C241 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=241655 $Y=21815 $dt=11
C242 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=241950 $Y=37085 $dt=11
C243 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=241950 $Y=48785 $dt=11
C244 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=241950 $Y=60485 $dt=11
C245 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=247695 $Y=10115 $dt=11
C246 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=247695 $Y=21815 $dt=11
C247 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=247990 $Y=37085 $dt=11
C248 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=247990 $Y=48785 $dt=11
C249 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=247990 $Y=60485 $dt=11
C250 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=253735 $Y=10115 $dt=11
C251 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=253735 $Y=21815 $dt=11
C252 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=254030 $Y=37085 $dt=11
C253 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=254030 $Y=48785 $dt=11
C254 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=254030 $Y=60485 $dt=11
C255 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=259775 $Y=10115 $dt=11
C256 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=259775 $Y=21815 $dt=11
C257 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=260070 $Y=37085 $dt=11
C258 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=260070 $Y=48785 $dt=11
C259 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=260070 $Y=60485 $dt=11
C260 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=265815 $Y=10115 $dt=11
C261 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=265815 $Y=21815 $dt=11
C262 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=266110 $Y=37085 $dt=11
C263 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=266110 $Y=48785 $dt=11
C264 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=266110 $Y=60485 $dt=11
C265 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=271855 $Y=10115 $dt=11
C266 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=271855 $Y=21815 $dt=11
C267 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=272150 $Y=37085 $dt=11
C268 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=272150 $Y=48785 $dt=11
C269 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=272150 $Y=60485 $dt=11
C270 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=277895 $Y=10115 $dt=11
C271 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=277895 $Y=21815 $dt=11
C272 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=278190 $Y=37085 $dt=11
C273 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=278190 $Y=48785 $dt=11
C274 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=278190 $Y=60485 $dt=11
C275 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=283935 $Y=10115 $dt=11
C276 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=283935 $Y=21815 $dt=11
C277 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=284230 $Y=37085 $dt=11
C278 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=284230 $Y=48785 $dt=11
C279 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=284230 $Y=60485 $dt=11
C280 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=289975 $Y=10115 $dt=11
C281 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=289975 $Y=21815 $dt=11
C282 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=290270 $Y=37085 $dt=11
C283 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=290270 $Y=48785 $dt=11
C284 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=290270 $Y=60485 $dt=11
C285 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=296015 $Y=10115 $dt=11
C286 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=296015 $Y=21815 $dt=11
C287 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=296310 $Y=37085 $dt=11
C288 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=296310 $Y=48785 $dt=11
C289 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=296310 $Y=60485 $dt=11
C290 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=302055 $Y=10115 $dt=11
C291 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=302055 $Y=21815 $dt=11
C292 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=302350 $Y=37085 $dt=11
C293 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=302350 $Y=48785 $dt=11
C294 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=302350 $Y=60485 $dt=11
C295 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=308095 $Y=10115 $dt=11
C296 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=308095 $Y=21815 $dt=11
C297 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=308390 $Y=37085 $dt=11
C298 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=308390 $Y=48785 $dt=11
C299 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=308390 $Y=60485 $dt=11
C300 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=314135 $Y=10115 $dt=11
C301 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=314135 $Y=21815 $dt=11
C302 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=314430 $Y=37085 $dt=11
C303 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=314430 $Y=48785 $dt=11
C304 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=314430 $Y=60485 $dt=11
C305 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=320175 $Y=10115 $dt=11
C306 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=320175 $Y=21815 $dt=11
C307 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=320470 $Y=37085 $dt=11
C308 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=320470 $Y=48785 $dt=11
C309 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=320470 $Y=60485 $dt=11
C310 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=326215 $Y=10115 $dt=11
C311 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=326215 $Y=21815 $dt=11
C312 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=326510 $Y=37085 $dt=11
C313 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=326510 $Y=48785 $dt=11
C314 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=326510 $Y=60485 $dt=11
C315 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=332255 $Y=10115 $dt=11
C316 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=332255 $Y=21815 $dt=11
C317 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=332550 $Y=37085 $dt=11
C318 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=332550 $Y=48785 $dt=11
C319 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=332550 $Y=60485 $dt=11
C320 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=338295 $Y=10115 $dt=11
C321 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=338295 $Y=21815 $dt=11
C322 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=338590 $Y=37085 $dt=11
C323 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=338590 $Y=48785 $dt=11
C324 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=338590 $Y=60485 $dt=11
C325 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=344335 $Y=10115 $dt=11
C326 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=344335 $Y=21815 $dt=11
C327 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=344630 $Y=37085 $dt=11
C328 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=344630 $Y=48785 $dt=11
C329 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=344630 $Y=60485 $dt=11
C330 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=350375 $Y=10115 $dt=11
C331 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=350375 $Y=21815 $dt=11
C332 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=350670 $Y=37085 $dt=11
C333 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=350670 $Y=48785 $dt=11
C334 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=350670 $Y=60485 $dt=11
C335 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=356415 $Y=10115 $dt=11
C336 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=356415 $Y=21815 $dt=11
C337 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=356710 $Y=37085 $dt=11
C338 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=356710 $Y=48785 $dt=11
C339 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=356710 $Y=60485 $dt=11
C340 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=362455 $Y=10115 $dt=11
C341 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=362455 $Y=21815 $dt=11
C342 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=362750 $Y=37085 $dt=11
C343 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=362750 $Y=48785 $dt=11
C344 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=362750 $Y=60485 $dt=11
C345 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=368495 $Y=10115 $dt=11
C346 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=368495 $Y=21815 $dt=11
C347 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=368790 $Y=37085 $dt=11
C348 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=368790 $Y=48785 $dt=11
C349 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=368790 $Y=60485 $dt=11
C350 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=374535 $Y=10115 $dt=11
C351 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=374535 $Y=21815 $dt=11
C352 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=374830 $Y=37085 $dt=11
C353 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=374830 $Y=48785 $dt=11
C354 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=374830 $Y=60485 $dt=11
C355 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=380575 $Y=10115 $dt=11
C356 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=380575 $Y=21815 $dt=11
C357 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=380870 $Y=37085 $dt=11
C358 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=380870 $Y=48785 $dt=11
C359 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=380870 $Y=60485 $dt=11
C360 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=386615 $Y=10115 $dt=11
C361 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=386615 $Y=21815 $dt=11
C362 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=386910 $Y=37085 $dt=11
C363 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=386910 $Y=48785 $dt=11
C364 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=386910 $Y=60485 $dt=11
C365 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=392655 $Y=10115 $dt=11
C366 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=392655 $Y=21815 $dt=11
C367 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=392950 $Y=37085 $dt=11
C368 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=392950 $Y=48785 $dt=11
C369 3 4 area=6.3936e-11 perimeter=3.372e-05 $[csf4a] $X=392950 $Y=60485 $dt=11
.ends MASCO__P2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724655180280                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724655180280 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724655180280

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724655180281                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724655180281 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724655180281

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724655180284                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724655180284 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724655180284

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_724655180285                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_724655180285 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_724655180285

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724655180287                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724655180287 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_724655180287

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724655180288                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724655180288 1 2
** N=2 EP=2 FDC=0
.ends VIA1_C_CDNS_724655180288

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_724655180289                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_724655180289 1 2
** N=2 EP=2 FDC=0
.ends VIA1_C_CDNS_724655180289

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246551802819                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246551802819 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246551802819

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7246551802821                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7246551802821 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7246551802821

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_7246551802822                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_7246551802822 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_7246551802822

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_7246551802823                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_7246551802823 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_7246551802823

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246551802824                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246551802824 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246551802824

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_7246551802825                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_7246551802825 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_7246551802825

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_7246551802826                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_7246551802826 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_7246551802826

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_7246551802827                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_7246551802827 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_7246551802827

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_7246551802829                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_7246551802829 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_7246551802829

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA3_C_CDNS_7246551802830                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA3_C_CDNS_7246551802830 1
** N=1 EP=1 FDC=0
.ends VIA3_C_CDNS_7246551802830

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246551802835                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246551802835 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246551802835

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246551802836                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246551802836 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246551802836

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246551802837                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246551802837 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246551802837

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246551802839                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246551802839 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246551802839

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246551802841                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246551802841 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246551802841

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIATP_C_CDNS_7246551802844                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIATP_C_CDNS_7246551802844 1
** N=1 EP=1 FDC=0
.ends VIATP_C_CDNS_7246551802844

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ped_CDNS_724655180281                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ped_CDNS_724655180281 1 2 3 4
** N=4 EP=4 FDC=12
X0 2 4 3 1 LDDP w=5e-05 l=9.4e-07 ad=2.19714e-10 pd=8.94366e-05 adio=4.2498e-10 pdio=2.57015e-05 extlay=1 $[ped] $X=-2270 $Y=0 $dt=1
X1 2 4 3 1 LDDP w=5e-05 l=9.4e-07 ad=2.19714e-10 pd=8.94366e-05 adio=4.2498e-10 pdio=2.57015e-05 extlay=1 $[ped] $X=6530 $Y=0 $dt=1
X2 2 4 3 1 LDDP w=5e-05 l=9.4e-07 ad=2.19714e-10 pd=8.94366e-05 adio=4.2498e-10 pdio=2.57015e-05 extlay=1 $[ped] $X=15330 $Y=0 $dt=1
X3 2 4 3 1 LDDP w=5e-05 l=9.4e-07 ad=2.19714e-10 pd=8.94366e-05 adio=4.2498e-10 pdio=2.57015e-05 extlay=1 $[ped] $X=24130 $Y=0 $dt=1
X4 2 4 3 1 LDDP w=5e-05 l=9.4e-07 ad=2.19714e-10 pd=8.94366e-05 adio=4.2498e-10 pdio=2.57015e-05 extlay=1 $[ped] $X=32930 $Y=0 $dt=1
X5 2 4 3 1 LDDP w=5e-05 l=9.4e-07 ad=2.19714e-10 pd=8.94366e-05 adio=4.2498e-10 pdio=2.57015e-05 extlay=1 $[ped] $X=41730 $Y=0 $dt=1
X6 2 4 3 1 LDDP w=5e-05 l=9.4e-07 ad=2.19714e-10 pd=8.94366e-05 adio=4.2498e-10 pdio=2.57015e-05 extlay=1 $[ped] $X=50530 $Y=0 $dt=1
X7 2 4 3 1 LDDP w=5e-05 l=9.4e-07 ad=2.19714e-10 pd=8.94366e-05 adio=4.2498e-10 pdio=2.57015e-05 extlay=1 $[ped] $X=59330 $Y=0 $dt=1
X8 2 4 3 1 LDDP w=5e-05 l=9.4e-07 ad=2.19714e-10 pd=8.94366e-05 adio=4.2498e-10 pdio=2.57015e-05 extlay=1 $[ped] $X=68130 $Y=0 $dt=1
X9 2 4 3 1 LDDP w=5e-05 l=9.4e-07 ad=2.19714e-10 pd=8.94366e-05 adio=4.2498e-10 pdio=2.57015e-05 extlay=1 $[ped] $X=76930 $Y=0 $dt=1
X10 2 4 3 1 LDDP w=5e-05 l=9.4e-07 ad=2.19714e-10 pd=8.94366e-05 adio=4.2498e-10 pdio=2.57015e-05 extlay=1 $[ped] $X=85730 $Y=0 $dt=1
X11 2 4 3 1 LDDP w=5e-05 l=9.4e-07 ad=2.19714e-10 pd=8.94366e-05 adio=4.2498e-10 pdio=2.57015e-05 extlay=1 $[ped] $X=94530 $Y=0 $dt=1
.ends ped_CDNS_724655180281

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nedia_CDNS_724655180282                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nedia_CDNS_724655180282 1 2 3 4
** N=4 EP=4 FDC=1
X0 2 4 3 1 LDDN w=2e-05 l=1.25e-06 adio=7.56916e-10 pdio=0.00010535 extlay=1 $[nedia] $X=-680 $Y=-4850 $dt=0
.ends nedia_CDNS_724655180282

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_724655180283                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_724655180283 1 2 3 4
** N=4 EP=4 FDC=1
M0 3 2 1 4 ne3 L=3.5e-07 W=2.2e-07 AD=1.984e-13 AS=1.984e-13 PD=1.88e-06 PS=1.88e-06 $X=0 $Y=0 $dt=2
.ends ne3_CDNS_724655180283

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_724655180285                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_724655180285 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.0002029 W=2e-06 $[rpp1k1_3] $SUB=3 $X=-2220 $Y=0 $dt=10
.ends rpp1k1_3_CDNS_724655180285

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: dsba_CDNS_724655180286                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt dsba_CDNS_724655180286 1 2 3
** N=623 EP=3 FDC=21
D0 1 2 p_dwhn AREA=6.69221e-10 PJ=0.00022132 perimeter=0.00022132 $X=-3330 $Y=-3970 $dt=6
D1 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=1390 $Y=1050 $dt=8
D2 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=5350 $Y=1050 $dt=8
D3 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=9310 $Y=1050 $dt=8
D4 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=13270 $Y=1050 $dt=8
D5 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=17230 $Y=1050 $dt=8
D6 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=21190 $Y=1050 $dt=8
D7 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=25150 $Y=1050 $dt=8
D8 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=29110 $Y=1050 $dt=8
D9 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=33070 $Y=1050 $dt=8
D10 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=37030 $Y=1050 $dt=8
D11 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=40990 $Y=1050 $dt=8
D12 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=44950 $Y=1050 $dt=8
D13 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=48910 $Y=1050 $dt=8
D14 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=52870 $Y=1050 $dt=8
D15 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=56830 $Y=1050 $dt=8
D16 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=60790 $Y=1050 $dt=8
D17 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=64750 $Y=1050 $dt=8
D18 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=68710 $Y=1050 $dt=8
D19 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=72670 $Y=1050 $dt=8
D20 3 2 dsba AREA=1.41e-11 PJ=3.188e-05 perimeter=3.188e-05 $SUB=1 $X=76630 $Y=1050 $dt=8
.ends dsba_CDNS_724655180286

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: dpp20_CDNS_724655180287                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt dpp20_CDNS_724655180287 1 2 3
** N=3 EP=3 FDC=2
D0 1 2 p_ddnw AREA=1.12107e-09 PJ=0.00016136 perimeter=0.00016136 $X=-6420 $Y=-6420 $dt=5
D1 3 2 dpp20 AREA=2.5e-10 PJ=0.00011 perimeter=0.00011 $X=0 $Y=0 $dt=7
.ends dpp20_CDNS_724655180287

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_724655180288                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_724655180288 1 2 3
** N=3 EP=3 FDC=1
R0 2 1 L=0.0002537 W=2e-06 $[rpp1k1_3] $SUB=3 $X=-2220 $Y=0 $dt=10
.ends rpp1k1_3_CDNS_724655180288

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_724655180289                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_724655180289 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
M0 3 2 1 1 pe3 L=3e-07 W=4.4e-07 AD=2.112e-13 AS=2.112e-13 PD=1.84e-06 PS=1.84e-06 $X=0 $Y=0 $dt=3
.ends pe3_CDNS_724655180289

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X11                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X11 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7246551802815 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7246551802815 $T=500 1500 0 0 $X=0 $Y=1000
X2 1 VIATP_C_CDNS_7246551802815 $T=500 2500 0 0 $X=0 $Y=2000
X3 1 VIATP_C_CDNS_7246551802815 $T=500 3500 0 0 $X=0 $Y=3000
X4 1 VIATP_C_CDNS_7246551802815 $T=500 4500 0 0 $X=0 $Y=4000
X5 1 VIATP_C_CDNS_7246551802815 $T=500 5500 0 0 $X=0 $Y=5000
X6 1 VIATP_C_CDNS_7246551802815 $T=500 6500 0 0 $X=0 $Y=6000
.ends MASCO__X11

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__X9                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__X9 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7246551802815 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7246551802815 $T=500 2500 0 0 $X=0 $Y=2000
X2 1 VIATP_C_CDNS_7246551802815 $T=500 4500 0 0 $X=0 $Y=4000
X3 1 VIATP_C_CDNS_7246551802815 $T=500 6500 0 0 $X=0 $Y=6000
X4 1 VIATP_C_CDNS_7246551802815 $T=500 8500 0 0 $X=0 $Y=8000
X5 1 VIATP_C_CDNS_7246551802815 $T=500 10500 0 0 $X=0 $Y=10000
X6 1 VIATP_C_CDNS_7246551802815 $T=500 12500 0 0 $X=0 $Y=12000
X7 1 VIATP_C_CDNS_7246551802815 $T=500 14500 0 0 $X=0 $Y=14000
X8 1 VIATP_C_CDNS_7246551802815 $T=500 16500 0 0 $X=0 $Y=16000
.ends MASCO__X9

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y13                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y13 1
** N=1 EP=1 FDC=0
X0 1 MASCO__X9 $T=0 0 0 0 $X=0 $Y=0
X1 1 MASCO__X9 $T=2000 0 0 0 $X=2000 $Y=0
X2 1 MASCO__X9 $T=4000 0 0 0 $X=4000 $Y=0
X3 1 MASCO__X9 $T=6000 0 0 0 $X=6000 $Y=0
.ends MASCO__Y13

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y14                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y14 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7246551802831 $T=500 750 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7246551802831 $T=1500 750 0 0 $X=1000 $Y=0
X2 1 VIATP_C_CDNS_7246551802831 $T=2500 750 0 0 $X=2000 $Y=0
X3 1 VIATP_C_CDNS_7246551802831 $T=3500 750 0 0 $X=3000 $Y=0
X4 1 VIATP_C_CDNS_7246551802831 $T=4500 750 0 0 $X=4000 $Y=0
X5 1 VIATP_C_CDNS_7246551802831 $T=5500 750 0 0 $X=5000 $Y=0
X6 1 VIATP_C_CDNS_7246551802831 $T=6500 750 0 0 $X=6000 $Y=0
X7 1 VIATP_C_CDNS_7246551802831 $T=7500 750 0 0 $X=7000 $Y=0
.ends MASCO__Y14

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y15                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y15 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7246551802815 $T=500 500 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7246551802815 $T=2500 500 0 0 $X=2000 $Y=0
X2 1 VIATP_C_CDNS_7246551802815 $T=4500 500 0 0 $X=4000 $Y=0
X3 1 VIATP_C_CDNS_7246551802815 $T=6500 500 0 0 $X=6000 $Y=0
.ends MASCO__Y15

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y16                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y16 1
** N=1 EP=1 FDC=0
X0 1 MASCO__X6 $T=0 0 0 0 $X=0 $Y=0
X1 1 MASCO__X6 $T=2000 0 0 0 $X=2000 $Y=0
X2 1 MASCO__X6 $T=4000 0 0 0 $X=4000 $Y=0
X3 1 MASCO__X6 $T=6000 0 0 0 $X=6000 $Y=0
.ends MASCO__Y16

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y17                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y17 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7246551802837 $T=500 440 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7246551802837 $T=1500 440 0 0 $X=1000 $Y=0
X2 1 VIATP_C_CDNS_7246551802837 $T=2500 440 0 0 $X=2000 $Y=0
X3 1 VIATP_C_CDNS_7246551802837 $T=3500 440 0 0 $X=3000 $Y=0
X4 1 VIATP_C_CDNS_7246551802837 $T=4500 440 0 0 $X=4000 $Y=0
X5 1 VIATP_C_CDNS_7246551802837 $T=5500 440 0 0 $X=5000 $Y=0
X6 1 VIATP_C_CDNS_7246551802837 $T=6500 440 0 0 $X=6000 $Y=0
X7 1 VIATP_C_CDNS_7246551802837 $T=7500 440 0 0 $X=7000 $Y=0
X8 1 VIATP_C_CDNS_7246551802837 $T=8500 440 0 0 $X=8000 $Y=0
X9 1 VIATP_C_CDNS_7246551802837 $T=9500 440 0 0 $X=9000 $Y=0
X10 1 VIATP_C_CDNS_7246551802837 $T=10500 440 0 0 $X=10000 $Y=0
X11 1 VIATP_C_CDNS_7246551802837 $T=11500 440 0 0 $X=11000 $Y=0
.ends MASCO__Y17

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y18                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y18 1
** N=1 EP=1 FDC=0
X0 1 VIATP_C_CDNS_7246551802833 $T=500 620 0 0 $X=0 $Y=0
X1 1 VIATP_C_CDNS_7246551802833 $T=1500 620 0 0 $X=1000 $Y=0
X2 1 VIATP_C_CDNS_7246551802833 $T=2500 620 0 0 $X=2000 $Y=0
X3 1 VIATP_C_CDNS_7246551802833 $T=3500 620 0 0 $X=3000 $Y=0
X4 1 VIATP_C_CDNS_7246551802833 $T=4500 620 0 0 $X=4000 $Y=0
X5 1 VIATP_C_CDNS_7246551802833 $T=5500 620 0 0 $X=5000 $Y=0
.ends MASCO__Y18

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__P3                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__P3 1 2 3 4 5 6 7 8 9 10
** N=15 EP=10 FDC=51
X0 11 VIA1_C_CDNS_724655180280 $T=21770 115795 0 0 $X=21280 $Y=115565
X1 12 VIA1_C_CDNS_724655180280 $T=25090 115795 0 0 $X=24600 $Y=115565
X2 13 VIA1_C_CDNS_724655180280 $T=28410 115795 0 0 $X=27920 $Y=115565
X3 6 VIA1_C_CDNS_724655180281 $T=20690 112655 0 0 $X=20460 $Y=112165
X4 6 VIA1_C_CDNS_724655180281 $T=20690 114845 0 0 $X=20460 $Y=114355
X5 11 VIA1_C_CDNS_724655180281 $T=21600 112085 0 0 $X=21370 $Y=111595
X6 7 VIA1_C_CDNS_724655180281 $T=24010 112645 0 0 $X=23780 $Y=112155
X7 7 VIA1_C_CDNS_724655180281 $T=24010 114845 0 0 $X=23780 $Y=114355
X8 12 VIA1_C_CDNS_724655180281 $T=24945 112075 0 0 $X=24715 $Y=111585
X9 12 VIA1_C_CDNS_724655180281 $T=27330 112645 0 0 $X=27100 $Y=112155
X10 12 VIA1_C_CDNS_724655180281 $T=27330 114845 0 0 $X=27100 $Y=114355
X11 13 VIA1_C_CDNS_724655180281 $T=28265 112075 0 0 $X=28035 $Y=111585
X12 2 VIA1_C_CDNS_724655180284 $T=13275 213850 0 0 $X=12525 $Y=212840
X13 3 VIA1_C_CDNS_724655180284 $T=17590 194950 0 0 $X=16840 $Y=193940
X14 4 VIA1_C_CDNS_724655180284 $T=19435 176670 0 0 $X=18685 $Y=175660
X15 14 VIA1_C_CDNS_724655180284 $T=53360 176670 0 0 $X=52610 $Y=175660
X16 2 VIA1_C_CDNS_724655180284 $T=59720 213460 0 0 $X=58970 $Y=212450
X17 13 VIA2_C_CDNS_724655180285 $T=28430 116695 0 0 $X=28200 $Y=115685
X18 11 VIA2_C_CDNS_724655180285 $T=31955 137810 0 0 $X=31725 $Y=136800
X19 11 VIA2_C_CDNS_724655180285 $T=31955 157230 0 0 $X=31725 $Y=156220
X20 13 VIA2_C_CDNS_724655180285 $T=71980 137810 0 0 $X=71750 $Y=136800
X21 13 VIA2_C_CDNS_724655180285 $T=71980 157230 0 0 $X=71750 $Y=156220
X22 4 VIA1_C_CDNS_724655180287 $T=121395 130205 0 0 $X=121165 $Y=121915
X23 4 VIA1_C_CDNS_724655180287 $T=125355 130205 0 0 $X=125125 $Y=121915
X24 4 VIA1_C_CDNS_724655180287 $T=129315 130205 0 0 $X=129085 $Y=121915
X25 4 VIA1_C_CDNS_724655180287 $T=133275 130205 0 0 $X=133045 $Y=121915
X26 4 VIA1_C_CDNS_724655180287 $T=137240 130205 0 0 $X=137010 $Y=121915
X27 4 VIA1_C_CDNS_724655180287 $T=141200 130205 0 0 $X=140970 $Y=121915
X28 4 VIA1_C_CDNS_724655180287 $T=145160 130205 0 0 $X=144930 $Y=121915
X29 4 VIA1_C_CDNS_724655180287 $T=149120 130205 0 0 $X=148890 $Y=121915
X30 4 VIA1_C_CDNS_724655180287 $T=153075 130205 0 0 $X=152845 $Y=121915
X31 4 VIA1_C_CDNS_724655180287 $T=157035 130205 0 0 $X=156805 $Y=121915
X32 4 VIA1_C_CDNS_724655180287 $T=160995 130205 0 0 $X=160765 $Y=121915
X33 4 VIA1_C_CDNS_724655180287 $T=164955 130205 0 0 $X=164725 $Y=121915
X34 4 VIA1_C_CDNS_724655180287 $T=168920 130205 0 0 $X=168690 $Y=121915
X35 4 VIA1_C_CDNS_724655180287 $T=172880 130205 0 0 $X=172650 $Y=121915
X36 4 VIA1_C_CDNS_724655180287 $T=176840 130205 0 0 $X=176610 $Y=121915
X37 4 VIA1_C_CDNS_724655180287 $T=180800 130205 0 0 $X=180570 $Y=121915
X38 4 VIA1_C_CDNS_724655180287 $T=184755 130205 0 0 $X=184525 $Y=121915
X39 4 VIA1_C_CDNS_724655180287 $T=188715 130205 0 0 $X=188485 $Y=121915
X40 4 VIA1_C_CDNS_724655180287 $T=192675 130205 0 0 $X=192445 $Y=121915
X41 4 VIA1_C_CDNS_724655180287 $T=196635 130205 0 0 $X=196405 $Y=121915
X42 2 1 VIA1_C_CDNS_724655180288 $T=139395 209375 0 0 $X=129025 $Y=208885
X43 2 1 VIA1_C_CDNS_724655180288 $T=216215 209630 0 0 $X=205845 $Y=209140
X44 9 1 VIA1_C_CDNS_724655180289 $T=138730 203470 0 0 $X=114200 $Y=201575
X45 9 1 VIA1_C_CDNS_724655180289 $T=216095 203470 0 0 $X=191565 $Y=201575
X46 2 VIATP_C_CDNS_7246551802819 $T=269935 210810 0 0 $X=269060 $Y=210310
X47 2 VIATP_C_CDNS_7246551802819 $T=269935 211810 0 0 $X=269060 $Y=211310
X48 2 VIATP_C_CDNS_7246551802819 $T=269935 212810 0 0 $X=269060 $Y=212310
X49 2 VIATP_C_CDNS_7246551802819 $T=269935 213810 0 0 $X=269060 $Y=213310
X50 2 VIATP_C_CDNS_7246551802819 $T=269935 214810 0 0 $X=269060 $Y=214310
X51 2 VIATP_C_CDNS_7246551802819 $T=269935 215810 0 0 $X=269060 $Y=215310
X52 2 VIATP_C_CDNS_7246551802819 $T=269935 216810 0 0 $X=269060 $Y=216310
X53 2 VIATP_C_CDNS_7246551802819 $T=269935 218810 0 0 $X=269060 $Y=218310
X54 2 VIATP_C_CDNS_7246551802819 $T=269935 219810 0 0 $X=269060 $Y=219310
X55 2 VIATP_C_CDNS_7246551802819 $T=269935 220810 0 0 $X=269060 $Y=220310
X56 2 VIATP_C_CDNS_7246551802819 $T=269935 221810 0 0 $X=269060 $Y=221310
X57 2 VIATP_C_CDNS_7246551802819 $T=269935 222810 0 0 $X=269060 $Y=222310
X58 2 VIATP_C_CDNS_7246551802819 $T=269935 223810 0 0 $X=269060 $Y=223310
X59 2 VIATP_C_CDNS_7246551802819 $T=269935 224810 0 0 $X=269060 $Y=224310
X60 2 VIATP_C_CDNS_7246551802819 $T=269935 225810 0 0 $X=269060 $Y=225310
X61 2 VIATP_C_CDNS_7246551802819 $T=269935 226810 0 0 $X=269060 $Y=226310
X62 2 VIATP_C_CDNS_7246551802819 $T=269935 227810 0 0 $X=269060 $Y=227310
X63 2 VIATP_C_CDNS_7246551802819 $T=269935 228810 0 0 $X=269060 $Y=228310
X64 2 VIATP_C_CDNS_7246551802819 $T=269935 229810 0 0 $X=269060 $Y=229310
X65 2 VIATP_C_CDNS_7246551802819 $T=269935 230810 0 0 $X=269060 $Y=230310
X66 2 VIATP_C_CDNS_7246551802819 $T=269935 231810 0 0 $X=269060 $Y=231310
X67 2 VIATP_C_CDNS_7246551802819 $T=269935 233810 0 0 $X=269060 $Y=233310
X68 2 VIATP_C_CDNS_7246551802819 $T=269935 234810 0 0 $X=269060 $Y=234310
X69 2 VIATP_C_CDNS_7246551802819 $T=269935 235810 0 0 $X=269060 $Y=235310
X70 2 VIATP_C_CDNS_7246551802819 $T=269935 236810 0 0 $X=269060 $Y=236310
X71 2 VIATP_C_CDNS_7246551802819 $T=404685 210810 0 0 $X=403810 $Y=210310
X72 2 VIATP_C_CDNS_7246551802819 $T=404685 211810 0 0 $X=403810 $Y=211310
X73 2 VIATP_C_CDNS_7246551802819 $T=404685 212810 0 0 $X=403810 $Y=212310
X74 2 VIATP_C_CDNS_7246551802819 $T=404685 213810 0 0 $X=403810 $Y=213310
X75 2 VIATP_C_CDNS_7246551802819 $T=404685 214810 0 0 $X=403810 $Y=214310
X76 2 VIATP_C_CDNS_7246551802819 $T=404685 215810 0 0 $X=403810 $Y=215310
X77 2 VIATP_C_CDNS_7246551802819 $T=404685 216810 0 0 $X=403810 $Y=216310
X78 2 VIATP_C_CDNS_7246551802819 $T=404685 217810 0 0 $X=403810 $Y=217310
X79 2 VIATP_C_CDNS_7246551802819 $T=404685 218810 0 0 $X=403810 $Y=218310
X80 2 VIATP_C_CDNS_7246551802819 $T=404685 219810 0 0 $X=403810 $Y=219310
X81 2 VIATP_C_CDNS_7246551802819 $T=404685 220810 0 0 $X=403810 $Y=220310
X82 2 VIATP_C_CDNS_7246551802819 $T=404685 221810 0 0 $X=403810 $Y=221310
X83 2 VIATP_C_CDNS_7246551802819 $T=404685 222810 0 0 $X=403810 $Y=222310
X84 2 VIATP_C_CDNS_7246551802819 $T=404685 223810 0 0 $X=403810 $Y=223310
X85 2 VIATP_C_CDNS_7246551802819 $T=404685 224810 0 0 $X=403810 $Y=224310
X86 2 VIATP_C_CDNS_7246551802819 $T=404685 225810 0 0 $X=403810 $Y=225310
X87 2 VIATP_C_CDNS_7246551802819 $T=404685 226810 0 0 $X=403810 $Y=226310
X88 2 VIATP_C_CDNS_7246551802819 $T=404685 227810 0 0 $X=403810 $Y=227310
X89 2 VIATP_C_CDNS_7246551802819 $T=404685 228810 0 0 $X=403810 $Y=228310
X90 2 VIATP_C_CDNS_7246551802819 $T=404685 229810 0 0 $X=403810 $Y=229310
X91 2 VIATP_C_CDNS_7246551802819 $T=404685 230810 0 0 $X=403810 $Y=230310
X92 2 VIATP_C_CDNS_7246551802819 $T=404685 231810 0 0 $X=403810 $Y=231310
X93 2 VIATP_C_CDNS_7246551802819 $T=404685 232810 0 0 $X=403810 $Y=232310
X94 2 VIATP_C_CDNS_7246551802819 $T=404685 233810 0 0 $X=403810 $Y=233310
X95 2 VIATP_C_CDNS_7246551802819 $T=404685 234810 0 0 $X=403810 $Y=234310
X96 2 VIATP_C_CDNS_7246551802819 $T=404685 235810 0 0 $X=403810 $Y=235310
X97 2 VIATP_C_CDNS_7246551802819 $T=404685 236810 0 0 $X=403810 $Y=236310
X98 6 VIA2_C_CDNS_7246551802821 $T=20690 113985 0 0 $X=20460 $Y=113495
X99 7 VIA2_C_CDNS_7246551802821 $T=24010 113060 0 0 $X=23780 $Y=112570
X100 9 VIA3_C_CDNS_7246551802822 $T=232755 165610 0 0 $X=232020 $Y=165110
X101 9 VIA3_C_CDNS_7246551802822 $T=232755 167610 0 0 $X=232020 $Y=167110
X102 9 VIA3_C_CDNS_7246551802822 $T=232755 169610 0 0 $X=232020 $Y=169110
X103 9 VIA3_C_CDNS_7246551802822 $T=232755 171610 0 0 $X=232020 $Y=171110
X104 9 VIA3_C_CDNS_7246551802823 $T=234995 164610 0 0 $X=234495 $Y=164110
X105 9 VIA3_C_CDNS_7246551802823 $T=234995 166610 0 0 $X=234495 $Y=166110
X106 9 VIA3_C_CDNS_7246551802823 $T=234995 168610 0 0 $X=234495 $Y=168110
X107 9 VIA3_C_CDNS_7246551802823 $T=234995 170610 0 0 $X=234495 $Y=170110
X108 9 VIA3_C_CDNS_7246551802823 $T=236995 164610 0 0 $X=236495 $Y=164110
X109 9 VIA3_C_CDNS_7246551802823 $T=236995 166610 0 0 $X=236495 $Y=166110
X110 9 VIA3_C_CDNS_7246551802823 $T=236995 168610 0 0 $X=236495 $Y=168110
X111 9 VIA3_C_CDNS_7246551802823 $T=236995 170610 0 0 $X=236495 $Y=170110
X112 9 VIA3_C_CDNS_7246551802823 $T=238995 164610 0 0 $X=238495 $Y=164110
X113 9 VIA3_C_CDNS_7246551802823 $T=238995 166610 0 0 $X=238495 $Y=166110
X114 9 VIA3_C_CDNS_7246551802823 $T=238995 168610 0 0 $X=238495 $Y=168110
X115 9 VIA3_C_CDNS_7246551802823 $T=238995 170610 0 0 $X=238495 $Y=170110
X116 9 VIA3_C_CDNS_7246551802823 $T=240995 164610 0 0 $X=240495 $Y=164110
X117 9 VIA3_C_CDNS_7246551802823 $T=240995 166610 0 0 $X=240495 $Y=166110
X118 9 VIA3_C_CDNS_7246551802823 $T=240995 168610 0 0 $X=240495 $Y=168110
X119 9 VIA3_C_CDNS_7246551802823 $T=240995 170610 0 0 $X=240495 $Y=170110
X120 2 VIATP_C_CDNS_7246551802824 $T=376065 210810 0 0 $X=375795 $Y=210310
X121 2 VIATP_C_CDNS_7246551802824 $T=376065 211810 0 0 $X=375795 $Y=211310
X122 2 VIATP_C_CDNS_7246551802824 $T=376065 212810 0 0 $X=375795 $Y=212310
X123 2 VIATP_C_CDNS_7246551802824 $T=376065 213810 0 0 $X=375795 $Y=213310
X124 2 VIATP_C_CDNS_7246551802824 $T=376065 214810 0 0 $X=375795 $Y=214310
X125 2 VIATP_C_CDNS_7246551802824 $T=376065 215810 0 0 $X=375795 $Y=215310
X126 2 VIATP_C_CDNS_7246551802824 $T=376065 216810 0 0 $X=375795 $Y=216310
X127 2 VIATP_C_CDNS_7246551802824 $T=376065 217810 0 0 $X=375795 $Y=217310
X128 2 VIATP_C_CDNS_7246551802824 $T=376065 218810 0 0 $X=375795 $Y=218310
X129 2 VIATP_C_CDNS_7246551802824 $T=376065 219810 0 0 $X=375795 $Y=219310
X130 2 VIATP_C_CDNS_7246551802824 $T=376065 220810 0 0 $X=375795 $Y=220310
X131 2 VIATP_C_CDNS_7246551802824 $T=376065 221810 0 0 $X=375795 $Y=221310
X132 2 VIATP_C_CDNS_7246551802824 $T=376065 222810 0 0 $X=375795 $Y=222310
X133 2 VIATP_C_CDNS_7246551802824 $T=376065 223810 0 0 $X=375795 $Y=223310
X134 2 VIATP_C_CDNS_7246551802824 $T=376065 224810 0 0 $X=375795 $Y=224310
X135 2 VIATP_C_CDNS_7246551802824 $T=376065 225810 0 0 $X=375795 $Y=225310
X136 2 VIATP_C_CDNS_7246551802824 $T=376065 226810 0 0 $X=375795 $Y=226310
X137 2 VIATP_C_CDNS_7246551802824 $T=376065 227810 0 0 $X=375795 $Y=227310
X138 2 VIATP_C_CDNS_7246551802824 $T=376065 228810 0 0 $X=375795 $Y=228310
X139 2 VIATP_C_CDNS_7246551802824 $T=376065 229810 0 0 $X=375795 $Y=229310
X140 2 VIATP_C_CDNS_7246551802824 $T=376065 230810 0 0 $X=375795 $Y=230310
X141 2 VIATP_C_CDNS_7246551802824 $T=376065 231810 0 0 $X=375795 $Y=231310
X142 2 VIATP_C_CDNS_7246551802824 $T=376065 232810 0 0 $X=375795 $Y=232310
X143 2 VIATP_C_CDNS_7246551802824 $T=376065 233810 0 0 $X=375795 $Y=233310
X144 2 VIATP_C_CDNS_7246551802824 $T=376065 234810 0 0 $X=375795 $Y=234310
X145 2 VIATP_C_CDNS_7246551802824 $T=376065 235810 0 0 $X=375795 $Y=235310
X146 2 VIATP_C_CDNS_7246551802824 $T=376065 236810 0 0 $X=375795 $Y=236310
X147 9 VIA3_C_CDNS_7246551802825 $T=232755 164610 0 0 $X=232020 $Y=164110
X148 9 VIA3_C_CDNS_7246551802825 $T=232755 166610 0 0 $X=232020 $Y=166110
X149 9 VIA3_C_CDNS_7246551802825 $T=232755 168610 0 0 $X=232020 $Y=168110
X150 9 VIA3_C_CDNS_7246551802825 $T=232755 170610 0 0 $X=232020 $Y=170110
X151 9 VIA3_C_CDNS_7246551802826 $T=233995 164610 0 0 $X=233495 $Y=164110
X152 9 VIA3_C_CDNS_7246551802826 $T=233995 166610 0 0 $X=233495 $Y=166110
X153 9 VIA3_C_CDNS_7246551802826 $T=233995 168610 0 0 $X=233495 $Y=168110
X154 9 VIA3_C_CDNS_7246551802826 $T=233995 170610 0 0 $X=233495 $Y=170110
X155 9 VIA3_C_CDNS_7246551802826 $T=235995 164610 0 0 $X=235495 $Y=164110
X156 9 VIA3_C_CDNS_7246551802826 $T=235995 166610 0 0 $X=235495 $Y=166110
X157 9 VIA3_C_CDNS_7246551802826 $T=235995 168610 0 0 $X=235495 $Y=168110
X158 9 VIA3_C_CDNS_7246551802826 $T=235995 170610 0 0 $X=235495 $Y=170110
X159 9 VIA3_C_CDNS_7246551802826 $T=237995 164610 0 0 $X=237495 $Y=164110
X160 9 VIA3_C_CDNS_7246551802826 $T=237995 166610 0 0 $X=237495 $Y=166110
X161 9 VIA3_C_CDNS_7246551802826 $T=237995 168610 0 0 $X=237495 $Y=168110
X162 9 VIA3_C_CDNS_7246551802826 $T=237995 170610 0 0 $X=237495 $Y=170110
X163 9 VIA3_C_CDNS_7246551802826 $T=239995 164610 0 0 $X=239495 $Y=164110
X164 9 VIA3_C_CDNS_7246551802826 $T=239995 166610 0 0 $X=239495 $Y=166110
X165 9 VIA3_C_CDNS_7246551802826 $T=239995 168610 0 0 $X=239495 $Y=168110
X166 9 VIA3_C_CDNS_7246551802826 $T=239995 170610 0 0 $X=239495 $Y=170110
X167 9 VIA3_C_CDNS_7246551802827 $T=234995 165610 0 0 $X=234495 $Y=165110
X168 9 VIA3_C_CDNS_7246551802827 $T=234995 167610 0 0 $X=234495 $Y=167110
X169 9 VIA3_C_CDNS_7246551802827 $T=234995 169610 0 0 $X=234495 $Y=169110
X170 9 VIA3_C_CDNS_7246551802827 $T=234995 171610 0 0 $X=234495 $Y=171110
X171 9 VIA3_C_CDNS_7246551802827 $T=236995 165610 0 0 $X=236495 $Y=165110
X172 9 VIA3_C_CDNS_7246551802827 $T=236995 167610 0 0 $X=236495 $Y=167110
X173 9 VIA3_C_CDNS_7246551802827 $T=236995 169610 0 0 $X=236495 $Y=169110
X174 9 VIA3_C_CDNS_7246551802827 $T=236995 171610 0 0 $X=236495 $Y=171110
X175 9 VIA3_C_CDNS_7246551802827 $T=238995 165610 0 0 $X=238495 $Y=165110
X176 9 VIA3_C_CDNS_7246551802827 $T=238995 167610 0 0 $X=238495 $Y=167110
X177 9 VIA3_C_CDNS_7246551802827 $T=238995 169610 0 0 $X=238495 $Y=169110
X178 9 VIA3_C_CDNS_7246551802827 $T=238995 171610 0 0 $X=238495 $Y=171110
X179 9 VIA3_C_CDNS_7246551802827 $T=240995 165610 0 0 $X=240495 $Y=165110
X180 9 VIA3_C_CDNS_7246551802827 $T=240995 167610 0 0 $X=240495 $Y=167110
X181 9 VIA3_C_CDNS_7246551802827 $T=240995 169610 0 0 $X=240495 $Y=169110
X182 9 VIA3_C_CDNS_7246551802827 $T=240995 171610 0 0 $X=240495 $Y=171110
X183 9 VIA3_C_CDNS_7246551802829 $T=233995 172860 0 0 $X=233495 $Y=172110
X184 9 VIA3_C_CDNS_7246551802829 $T=235995 172860 0 0 $X=235495 $Y=172110
X185 9 VIA3_C_CDNS_7246551802829 $T=237995 172860 0 0 $X=237495 $Y=172110
X186 9 VIA3_C_CDNS_7246551802829 $T=239995 172860 0 0 $X=239495 $Y=172110
X187 9 VIA3_C_CDNS_7246551802830 $T=234995 172860 0 0 $X=234495 $Y=172110
X188 9 VIA3_C_CDNS_7246551802830 $T=236995 172860 0 0 $X=236495 $Y=172110
X189 9 VIA3_C_CDNS_7246551802830 $T=238995 172860 0 0 $X=238495 $Y=172110
X190 9 VIA3_C_CDNS_7246551802830 $T=240995 172860 0 0 $X=240495 $Y=172110
X191 2 VIATP_C_CDNS_7246551802831 $T=377310 238060 0 0 $X=376810 $Y=237310
X192 2 VIATP_C_CDNS_7246551802831 $T=378310 238060 0 0 $X=377810 $Y=237310
X193 2 VIATP_C_CDNS_7246551802831 $T=379310 238060 0 0 $X=378810 $Y=237310
X194 2 VIATP_C_CDNS_7246551802831 $T=380310 238060 0 0 $X=379810 $Y=237310
X195 2 VIATP_C_CDNS_7246551802831 $T=381310 238060 0 0 $X=380810 $Y=237310
X196 2 VIATP_C_CDNS_7246551802831 $T=382310 238060 0 0 $X=381810 $Y=237310
X197 2 VIATP_C_CDNS_7246551802831 $T=383310 238060 0 0 $X=382810 $Y=237310
X198 2 VIATP_C_CDNS_7246551802831 $T=384310 238060 0 0 $X=383810 $Y=237310
X199 2 VIATP_C_CDNS_7246551802831 $T=385310 238060 0 0 $X=384810 $Y=237310
X200 2 VIATP_C_CDNS_7246551802831 $T=386310 238060 0 0 $X=385810 $Y=237310
X201 2 VIATP_C_CDNS_7246551802831 $T=387310 238060 0 0 $X=386810 $Y=237310
X202 2 VIATP_C_CDNS_7246551802831 $T=388310 238060 0 0 $X=387810 $Y=237310
X203 2 VIATP_C_CDNS_7246551802831 $T=389310 238060 0 0 $X=388810 $Y=237310
X204 2 VIATP_C_CDNS_7246551802831 $T=390310 238060 0 0 $X=389810 $Y=237310
X205 2 VIATP_C_CDNS_7246551802831 $T=391310 238060 0 0 $X=390810 $Y=237310
X206 2 VIATP_C_CDNS_7246551802831 $T=392310 238060 0 0 $X=391810 $Y=237310
X207 2 VIATP_C_CDNS_7246551802831 $T=393310 238060 0 0 $X=392810 $Y=237310
X208 2 VIATP_C_CDNS_7246551802831 $T=394310 238060 0 0 $X=393810 $Y=237310
X209 2 VIATP_C_CDNS_7246551802831 $T=395310 238060 0 0 $X=394810 $Y=237310
X210 2 VIATP_C_CDNS_7246551802831 $T=396310 238060 0 0 $X=395810 $Y=237310
X211 2 VIATP_C_CDNS_7246551802831 $T=397310 238060 0 0 $X=396810 $Y=237310
X212 2 VIATP_C_CDNS_7246551802831 $T=398310 238060 0 0 $X=397810 $Y=237310
X213 2 VIATP_C_CDNS_7246551802831 $T=399310 238060 0 0 $X=398810 $Y=237310
X214 2 VIATP_C_CDNS_7246551802831 $T=400310 238060 0 0 $X=399810 $Y=237310
X215 2 VIATP_C_CDNS_7246551802831 $T=401310 238060 0 0 $X=400810 $Y=237310
X216 2 VIATP_C_CDNS_7246551802831 $T=402310 238060 0 0 $X=401810 $Y=237310
X217 2 VIATP_C_CDNS_7246551802831 $T=403310 238060 0 0 $X=402810 $Y=237310
X218 9 VIATP_C_CDNS_7246551802833 $T=257995 172730 0 0 $X=257495 $Y=172110
X219 9 VIATP_C_CDNS_7246551802833 $T=258995 172730 0 0 $X=258495 $Y=172110
X220 9 VIATP_C_CDNS_7246551802833 $T=259995 172730 0 0 $X=259495 $Y=172110
X221 9 VIATP_C_CDNS_7246551802833 $T=260995 172730 0 0 $X=260495 $Y=172110
X222 9 VIATP_C_CDNS_7246551802833 $T=261995 172730 0 0 $X=261495 $Y=172110
X223 9 VIATP_C_CDNS_7246551802833 $T=262995 172730 0 0 $X=262495 $Y=172110
X224 9 VIATP_C_CDNS_7246551802833 $T=263995 172730 0 0 $X=263495 $Y=172110
X225 9 VIATP_C_CDNS_7246551802833 $T=264995 172730 0 0 $X=264495 $Y=172110
X226 9 VIATP_C_CDNS_7246551802833 $T=265995 172730 0 0 $X=265495 $Y=172110
X227 9 VIATP_C_CDNS_7246551802833 $T=266995 172730 0 0 $X=266495 $Y=172110
X228 9 VIATP_C_CDNS_7246551802833 $T=365995 172730 0 0 $X=365495 $Y=172110
X229 9 VIATP_C_CDNS_7246551802833 $T=366995 172730 0 0 $X=366495 $Y=172110
X230 9 VIATP_C_CDNS_7246551802833 $T=367995 172730 0 0 $X=367495 $Y=172110
X231 9 VIATP_C_CDNS_7246551802833 $T=368995 172730 0 0 $X=368495 $Y=172110
X232 9 VIATP_C_CDNS_7246551802833 $T=369995 172730 0 0 $X=369495 $Y=172110
X233 9 VIATP_C_CDNS_7246551802833 $T=370995 172730 0 0 $X=370495 $Y=172110
X234 9 VIATP_C_CDNS_7246551802833 $T=371995 172730 0 0 $X=371495 $Y=172110
X235 9 VIATP_C_CDNS_7246551802833 $T=372995 172730 0 0 $X=372495 $Y=172110
X236 9 VIATP_C_CDNS_7246551802833 $T=373995 172730 0 0 $X=373495 $Y=172110
X237 2 VIATP_C_CDNS_7246551802833 $T=374310 209690 0 0 $X=373810 $Y=209070
X238 9 VIATP_C_CDNS_7246551802833 $T=374995 172730 0 0 $X=374495 $Y=172110
X239 2 VIATP_C_CDNS_7246551802833 $T=375310 209690 0 0 $X=374810 $Y=209070
X240 2 VIATP_C_CDNS_7246551802833 $T=377310 209690 0 0 $X=376810 $Y=209070
X241 9 VIATP_C_CDNS_7246551802833 $T=377995 172730 0 0 $X=377495 $Y=172110
X242 2 VIATP_C_CDNS_7246551802833 $T=378310 209690 0 0 $X=377810 $Y=209070
X243 9 VIATP_C_CDNS_7246551802833 $T=378995 172730 0 0 $X=378495 $Y=172110
X244 2 VIATP_C_CDNS_7246551802833 $T=379310 209690 0 0 $X=378810 $Y=209070
X245 9 VIATP_C_CDNS_7246551802833 $T=379995 172730 0 0 $X=379495 $Y=172110
X246 2 VIATP_C_CDNS_7246551802833 $T=380310 209690 0 0 $X=379810 $Y=209070
X247 9 VIATP_C_CDNS_7246551802833 $T=380995 172730 0 0 $X=380495 $Y=172110
X248 2 VIATP_C_CDNS_7246551802833 $T=381310 209690 0 0 $X=380810 $Y=209070
X249 9 VIATP_C_CDNS_7246551802833 $T=381995 172730 0 0 $X=381495 $Y=172110
X250 2 VIATP_C_CDNS_7246551802833 $T=382310 209690 0 0 $X=381810 $Y=209070
X251 9 VIATP_C_CDNS_7246551802833 $T=382995 172730 0 0 $X=382495 $Y=172110
X252 2 VIATP_C_CDNS_7246551802833 $T=383310 209690 0 0 $X=382810 $Y=209070
X253 9 VIATP_C_CDNS_7246551802833 $T=383995 172730 0 0 $X=383495 $Y=172110
X254 2 VIATP_C_CDNS_7246551802833 $T=384310 209690 0 0 $X=383810 $Y=209070
X255 9 VIATP_C_CDNS_7246551802833 $T=384995 172730 0 0 $X=384495 $Y=172110
X256 2 VIATP_C_CDNS_7246551802833 $T=385310 209690 0 0 $X=384810 $Y=209070
X257 9 VIATP_C_CDNS_7246551802833 $T=385995 144490 0 0 $X=385495 $Y=143870
X258 9 VIATP_C_CDNS_7246551802833 $T=385995 172730 0 0 $X=385495 $Y=172110
X259 2 VIATP_C_CDNS_7246551802833 $T=386310 209690 0 0 $X=385810 $Y=209070
X260 9 VIATP_C_CDNS_7246551802833 $T=386995 144490 0 0 $X=386495 $Y=143870
X261 9 VIATP_C_CDNS_7246551802833 $T=386995 172730 0 0 $X=386495 $Y=172110
X262 2 VIATP_C_CDNS_7246551802833 $T=387310 209690 0 0 $X=386810 $Y=209070
X263 9 VIATP_C_CDNS_7246551802833 $T=387995 144490 0 0 $X=387495 $Y=143870
X264 9 VIATP_C_CDNS_7246551802833 $T=387995 172730 0 0 $X=387495 $Y=172110
X265 2 VIATP_C_CDNS_7246551802833 $T=388310 209690 0 0 $X=387810 $Y=209070
X266 9 VIATP_C_CDNS_7246551802833 $T=388995 144490 0 0 $X=388495 $Y=143870
X267 9 VIATP_C_CDNS_7246551802833 $T=388995 172730 0 0 $X=388495 $Y=172110
X268 2 VIATP_C_CDNS_7246551802833 $T=389310 209690 0 0 $X=388810 $Y=209070
X269 9 VIATP_C_CDNS_7246551802833 $T=389995 144490 0 0 $X=389495 $Y=143870
X270 9 VIATP_C_CDNS_7246551802833 $T=389995 172730 0 0 $X=389495 $Y=172110
X271 2 VIATP_C_CDNS_7246551802833 $T=390310 209690 0 0 $X=389810 $Y=209070
X272 9 VIATP_C_CDNS_7246551802833 $T=390995 144490 0 0 $X=390495 $Y=143870
X273 9 VIATP_C_CDNS_7246551802833 $T=390995 172730 0 0 $X=390495 $Y=172110
X274 2 VIATP_C_CDNS_7246551802833 $T=391310 209690 0 0 $X=390810 $Y=209070
X275 9 VIATP_C_CDNS_7246551802833 $T=391995 144490 0 0 $X=391495 $Y=143870
X276 9 VIATP_C_CDNS_7246551802833 $T=391995 172730 0 0 $X=391495 $Y=172110
X277 2 VIATP_C_CDNS_7246551802833 $T=392310 209690 0 0 $X=391810 $Y=209070
X278 9 VIATP_C_CDNS_7246551802833 $T=392995 144490 0 0 $X=392495 $Y=143870
X279 9 VIATP_C_CDNS_7246551802833 $T=392995 172730 0 0 $X=392495 $Y=172110
X280 2 VIATP_C_CDNS_7246551802833 $T=393310 209690 0 0 $X=392810 $Y=209070
X281 9 VIATP_C_CDNS_7246551802833 $T=393995 144490 0 0 $X=393495 $Y=143870
X282 9 VIATP_C_CDNS_7246551802833 $T=393995 172730 0 0 $X=393495 $Y=172110
X283 2 VIATP_C_CDNS_7246551802833 $T=394310 209690 0 0 $X=393810 $Y=209070
X284 9 VIATP_C_CDNS_7246551802833 $T=394995 144490 0 0 $X=394495 $Y=143870
X285 9 VIATP_C_CDNS_7246551802833 $T=394995 172730 0 0 $X=394495 $Y=172110
X286 2 VIATP_C_CDNS_7246551802833 $T=395310 209690 0 0 $X=394810 $Y=209070
X287 9 VIATP_C_CDNS_7246551802833 $T=395995 144490 0 0 $X=395495 $Y=143870
X288 9 VIATP_C_CDNS_7246551802833 $T=395995 172730 0 0 $X=395495 $Y=172110
X289 2 VIATP_C_CDNS_7246551802833 $T=396310 209690 0 0 $X=395810 $Y=209070
X290 9 VIATP_C_CDNS_7246551802833 $T=396995 144490 0 0 $X=396495 $Y=143870
X291 9 VIATP_C_CDNS_7246551802833 $T=396995 172730 0 0 $X=396495 $Y=172110
X292 2 VIATP_C_CDNS_7246551802833 $T=397310 209690 0 0 $X=396810 $Y=209070
X293 9 VIATP_C_CDNS_7246551802833 $T=397995 144490 0 0 $X=397495 $Y=143870
X294 9 VIATP_C_CDNS_7246551802833 $T=397995 172730 0 0 $X=397495 $Y=172110
X295 2 VIATP_C_CDNS_7246551802833 $T=398310 209690 0 0 $X=397810 $Y=209070
X296 9 VIATP_C_CDNS_7246551802833 $T=398995 144490 0 0 $X=398495 $Y=143870
X297 9 VIATP_C_CDNS_7246551802833 $T=398995 172730 0 0 $X=398495 $Y=172110
X298 2 VIATP_C_CDNS_7246551802833 $T=399310 209690 0 0 $X=398810 $Y=209070
X299 9 VIATP_C_CDNS_7246551802833 $T=399995 144490 0 0 $X=399495 $Y=143870
X300 9 VIATP_C_CDNS_7246551802833 $T=399995 172730 0 0 $X=399495 $Y=172110
X301 2 VIATP_C_CDNS_7246551802833 $T=400310 209690 0 0 $X=399810 $Y=209070
X302 9 VIATP_C_CDNS_7246551802833 $T=400995 144490 0 0 $X=400495 $Y=143870
X303 9 VIATP_C_CDNS_7246551802833 $T=400995 172730 0 0 $X=400495 $Y=172110
X304 2 VIATP_C_CDNS_7246551802833 $T=401310 209690 0 0 $X=400810 $Y=209070
X305 9 VIATP_C_CDNS_7246551802833 $T=401995 144490 0 0 $X=401495 $Y=143870
X306 9 VIATP_C_CDNS_7246551802833 $T=401995 172730 0 0 $X=401495 $Y=172110
X307 2 VIATP_C_CDNS_7246551802833 $T=402310 209690 0 0 $X=401810 $Y=209070
X308 9 VIATP_C_CDNS_7246551802833 $T=402995 144490 0 0 $X=402495 $Y=143870
X309 9 VIATP_C_CDNS_7246551802833 $T=402995 172730 0 0 $X=402495 $Y=172110
X310 2 VIATP_C_CDNS_7246551802833 $T=403310 209690 0 0 $X=402810 $Y=209070
X311 9 VIATP_C_CDNS_7246551802833 $T=403995 144490 0 0 $X=403495 $Y=143870
X312 9 VIATP_C_CDNS_7246551802833 $T=403995 172730 0 0 $X=403495 $Y=172110
X313 2 VIATP_C_CDNS_7246551802834 $T=373365 209690 0 0 $X=372925 $Y=209070
X314 2 VIATP_C_CDNS_7246551802835 $T=269935 209690 0 0 $X=269060 $Y=209070
X315 2 VIATP_C_CDNS_7246551802835 $T=404685 209690 0 0 $X=403810 $Y=209070
X316 2 VIATP_C_CDNS_7246551802836 $T=269935 238060 0 0 $X=269060 $Y=237310
X317 2 VIATP_C_CDNS_7246551802836 $T=404685 238060 0 0 $X=403810 $Y=237310
X318 2 VIATP_C_CDNS_7246551802837 $T=367310 217750 0 0 $X=366810 $Y=217310
X319 2 VIATP_C_CDNS_7246551802837 $T=368310 217750 0 0 $X=367810 $Y=217310
X320 2 VIATP_C_CDNS_7246551802837 $T=369310 217750 0 0 $X=368810 $Y=217310
X321 2 VIATP_C_CDNS_7246551802837 $T=370310 217750 0 0 $X=369810 $Y=217310
X322 2 VIATP_C_CDNS_7246551802837 $T=371310 217750 0 0 $X=370810 $Y=217310
X323 2 VIATP_C_CDNS_7246551802837 $T=372310 217750 0 0 $X=371810 $Y=217310
X324 2 VIATP_C_CDNS_7246551802837 $T=373310 217750 0 0 $X=372810 $Y=217310
X325 2 VIATP_C_CDNS_7246551802839 $T=259815 218810 0 0 $X=250570 $Y=218310
X326 2 VIATP_C_CDNS_7246551802839 $T=259815 219810 0 0 $X=250570 $Y=219310
X327 2 VIATP_C_CDNS_7246551802839 $T=259815 220810 0 0 $X=250570 $Y=220310
X328 2 VIATP_C_CDNS_7246551802839 $T=259815 221810 0 0 $X=250570 $Y=221310
X329 2 VIATP_C_CDNS_7246551802839 $T=259815 222810 0 0 $X=250570 $Y=222310
X330 2 VIATP_C_CDNS_7246551802839 $T=259815 223810 0 0 $X=250570 $Y=223310
X331 2 VIATP_C_CDNS_7246551802839 $T=259815 224810 0 0 $X=250570 $Y=224310
X332 2 VIATP_C_CDNS_7246551802839 $T=259815 225810 0 0 $X=250570 $Y=225310
X333 2 VIATP_C_CDNS_7246551802839 $T=259815 226810 0 0 $X=250570 $Y=226310
X334 2 VIATP_C_CDNS_7246551802839 $T=259815 227810 0 0 $X=250570 $Y=227310
X335 2 VIATP_C_CDNS_7246551802839 $T=259815 228810 0 0 $X=250570 $Y=228310
X336 2 VIATP_C_CDNS_7246551802839 $T=259815 229810 0 0 $X=250570 $Y=229310
X337 2 VIATP_C_CDNS_7246551802839 $T=259815 230810 0 0 $X=250570 $Y=230310
X338 2 VIATP_C_CDNS_7246551802839 $T=259815 231810 0 0 $X=250570 $Y=231310
X339 9 VIATP_C_CDNS_7246551802841 $T=405235 145610 0 0 $X=404495 $Y=145110
X340 9 VIATP_C_CDNS_7246551802841 $T=405235 146610 0 0 $X=404495 $Y=146110
X341 9 VIATP_C_CDNS_7246551802841 $T=405235 147610 0 0 $X=404495 $Y=147110
X342 9 VIATP_C_CDNS_7246551802841 $T=405235 148610 0 0 $X=404495 $Y=148110
X343 9 VIATP_C_CDNS_7246551802841 $T=405235 149610 0 0 $X=404495 $Y=149110
X344 9 VIATP_C_CDNS_7246551802841 $T=405235 150610 0 0 $X=404495 $Y=150110
X345 9 VIATP_C_CDNS_7246551802841 $T=405235 151610 0 0 $X=404495 $Y=151110
X346 9 VIATP_C_CDNS_7246551802841 $T=405235 152610 0 0 $X=404495 $Y=152110
X347 9 VIATP_C_CDNS_7246551802841 $T=405235 153610 0 0 $X=404495 $Y=153110
X348 9 VIATP_C_CDNS_7246551802841 $T=405235 154610 0 0 $X=404495 $Y=154110
X349 9 VIATP_C_CDNS_7246551802841 $T=405235 155610 0 0 $X=404495 $Y=155110
X350 9 VIATP_C_CDNS_7246551802841 $T=405235 156610 0 0 $X=404495 $Y=156110
X351 9 VIATP_C_CDNS_7246551802841 $T=405235 157610 0 0 $X=404495 $Y=157110
X352 9 VIATP_C_CDNS_7246551802841 $T=405235 158610 0 0 $X=404495 $Y=158110
X353 9 VIATP_C_CDNS_7246551802841 $T=405235 159610 0 0 $X=404495 $Y=159110
X354 9 VIATP_C_CDNS_7246551802841 $T=405235 160610 0 0 $X=404495 $Y=160110
X355 9 VIATP_C_CDNS_7246551802841 $T=405235 161610 0 0 $X=404495 $Y=161110
X356 9 VIATP_C_CDNS_7246551802841 $T=405235 162610 0 0 $X=404495 $Y=162110
X357 9 VIATP_C_CDNS_7246551802841 $T=405235 163610 0 0 $X=404495 $Y=163110
X358 9 VIATP_C_CDNS_7246551802841 $T=405235 164610 0 0 $X=404495 $Y=164110
X359 9 VIATP_C_CDNS_7246551802841 $T=405235 165610 0 0 $X=404495 $Y=165110
X360 9 VIATP_C_CDNS_7246551802841 $T=405235 166610 0 0 $X=404495 $Y=166110
X361 9 VIATP_C_CDNS_7246551802841 $T=405235 167610 0 0 $X=404495 $Y=167110
X362 9 VIATP_C_CDNS_7246551802841 $T=405235 168610 0 0 $X=404495 $Y=168110
X363 9 VIATP_C_CDNS_7246551802841 $T=405235 169610 0 0 $X=404495 $Y=169110
X364 9 VIATP_C_CDNS_7246551802841 $T=405235 170610 0 0 $X=404495 $Y=170110
X365 9 VIATP_C_CDNS_7246551802841 $T=405235 171610 0 0 $X=404495 $Y=171110
X366 9 VIATP_C_CDNS_7246551802842 $T=376745 155610 0 0 $X=376475 $Y=155110
X367 9 VIATP_C_CDNS_7246551802842 $T=376745 156610 0 0 $X=376475 $Y=156110
X368 9 VIATP_C_CDNS_7246551802842 $T=376745 157610 0 0 $X=376475 $Y=157110
X369 9 VIATP_C_CDNS_7246551802842 $T=376745 158610 0 0 $X=376475 $Y=158110
X370 9 VIATP_C_CDNS_7246551802842 $T=376745 159610 0 0 $X=376475 $Y=159110
X371 9 VIATP_C_CDNS_7246551802842 $T=376745 160610 0 0 $X=376475 $Y=160110
X372 9 VIATP_C_CDNS_7246551802842 $T=376745 161610 0 0 $X=376475 $Y=161110
X373 9 VIATP_C_CDNS_7246551802842 $T=376745 162610 0 0 $X=376475 $Y=162110
X374 9 VIATP_C_CDNS_7246551802842 $T=376745 163610 0 0 $X=376475 $Y=163110
X375 9 VIATP_C_CDNS_7246551802842 $T=376745 164610 0 0 $X=376475 $Y=164110
X376 9 VIATP_C_CDNS_7246551802842 $T=376745 165610 0 0 $X=376475 $Y=165110
X377 9 VIATP_C_CDNS_7246551802842 $T=376745 166610 0 0 $X=376475 $Y=166110
X378 9 VIATP_C_CDNS_7246551802842 $T=376745 167610 0 0 $X=376475 $Y=167110
X379 9 VIATP_C_CDNS_7246551802842 $T=376745 168610 0 0 $X=376475 $Y=168110
X380 9 VIATP_C_CDNS_7246551802842 $T=376745 169610 0 0 $X=376475 $Y=169110
X381 9 VIATP_C_CDNS_7246551802842 $T=376745 170610 0 0 $X=376475 $Y=170110
X382 9 VIATP_C_CDNS_7246551802842 $T=376745 171610 0 0 $X=376475 $Y=171110
X383 9 VIATP_C_CDNS_7246551802844 $T=405235 144490 0 0 $X=404495 $Y=143870
X384 9 VIATP_C_CDNS_7246551802844 $T=405235 172730 0 0 $X=404495 $Y=172110
X385 9 VIATP_C_CDNS_7246551802846 $T=232755 172730 0 0 $X=232025 $Y=172110
X386 9 VIATP_C_CDNS_7246551802847 $T=268645 155610 0 0 $X=268375 $Y=155110
X387 9 VIATP_C_CDNS_7246551802847 $T=268645 156610 0 0 $X=268375 $Y=156110
X388 9 VIATP_C_CDNS_7246551802847 $T=268645 157610 0 0 $X=268375 $Y=157110
X389 9 VIATP_C_CDNS_7246551802847 $T=268645 158610 0 0 $X=268375 $Y=158110
X390 9 VIATP_C_CDNS_7246551802847 $T=268645 159610 0 0 $X=268375 $Y=159110
X391 9 VIATP_C_CDNS_7246551802847 $T=268645 160610 0 0 $X=268375 $Y=160110
X392 9 VIATP_C_CDNS_7246551802847 $T=268645 161610 0 0 $X=268375 $Y=161110
X393 9 VIATP_C_CDNS_7246551802847 $T=268645 162610 0 0 $X=268375 $Y=162110
X394 9 VIATP_C_CDNS_7246551802847 $T=268645 163610 0 0 $X=268375 $Y=163110
X395 9 VIATP_C_CDNS_7246551802847 $T=268645 164610 0 0 $X=268375 $Y=164110
X396 9 VIATP_C_CDNS_7246551802847 $T=268645 165610 0 0 $X=268375 $Y=165110
X397 9 VIATP_C_CDNS_7246551802847 $T=268645 166610 0 0 $X=268375 $Y=166110
X398 9 VIATP_C_CDNS_7246551802847 $T=268645 167610 0 0 $X=268375 $Y=167110
X399 9 VIATP_C_CDNS_7246551802847 $T=268645 168610 0 0 $X=268375 $Y=168110
X400 9 VIATP_C_CDNS_7246551802847 $T=268645 169610 0 0 $X=268375 $Y=169110
X401 9 VIATP_C_CDNS_7246551802847 $T=268645 170610 0 0 $X=268375 $Y=170110
X402 9 VIATP_C_CDNS_7246551802847 $T=268645 171610 0 0 $X=268375 $Y=171110
X403 9 VIATP_C_CDNS_7246551802848 $T=232755 155610 0 0 $X=232025 $Y=155110
X404 9 VIATP_C_CDNS_7246551802848 $T=232755 156610 0 0 $X=232025 $Y=156110
X405 9 VIATP_C_CDNS_7246551802848 $T=232755 157610 0 0 $X=232025 $Y=157110
X406 9 VIATP_C_CDNS_7246551802848 $T=232755 158610 0 0 $X=232025 $Y=158110
X407 9 VIATP_C_CDNS_7246551802848 $T=232755 159610 0 0 $X=232025 $Y=159110
X408 9 VIATP_C_CDNS_7246551802848 $T=232755 160610 0 0 $X=232025 $Y=160110
X409 9 VIATP_C_CDNS_7246551802848 $T=232755 161610 0 0 $X=232025 $Y=161110
X410 9 VIATP_C_CDNS_7246551802848 $T=232755 162610 0 0 $X=232025 $Y=162110
X411 9 VIATP_C_CDNS_7246551802848 $T=232755 163610 0 0 $X=232025 $Y=163110
X412 9 VIATP_C_CDNS_7246551802848 $T=232755 164610 0 0 $X=232025 $Y=164110
X413 9 VIATP_C_CDNS_7246551802848 $T=232755 165610 0 0 $X=232025 $Y=165110
X414 9 VIATP_C_CDNS_7246551802848 $T=232755 166610 0 0 $X=232025 $Y=166110
X415 9 VIATP_C_CDNS_7246551802848 $T=232755 167610 0 0 $X=232025 $Y=167110
X416 9 VIATP_C_CDNS_7246551802848 $T=232755 168610 0 0 $X=232025 $Y=168110
X417 9 VIATP_C_CDNS_7246551802848 $T=232755 169610 0 0 $X=232025 $Y=169110
X418 9 VIATP_C_CDNS_7246551802848 $T=232755 170610 0 0 $X=232025 $Y=170110
X419 9 VIATP_C_CDNS_7246551802848 $T=232755 171610 0 0 $X=232025 $Y=171110
X420 1 9 2 15 ped_CDNS_724655180281 $T=370960 203710 0 180 $X=259210 $Y=163760
X421 1 3 4 11 nedia_CDNS_724655180282 $T=31955 142520 0 0 $X=15735 $Y=123130
X422 1 14 4 13 nedia_CDNS_724655180282 $T=71980 142520 0 0 $X=55760 $Y=123130
X423 8 6 11 1 ne3_CDNS_724655180283 $T=20540 111655 0 0 $X=19700 $Y=111235
X424 8 7 12 1 ne3_CDNS_724655180283 $T=23885 111645 0 0 $X=23045 $Y=111225
X425 8 12 13 1 ne3_CDNS_724655180283 $T=27205 111645 0 0 $X=26365 $Y=111225
X426 3 4 1 rpp1k1_3_CDNS_724655180285 $T=22985 175685 0 0 $X=19825 $Y=175465
X427 2 15 1 rpp1k1_3_CDNS_724655180285 $T=63010 196610 0 0 $X=59850 $Y=196390
X428 1 3 4 dsba_CDNS_724655180286 $T=119535 121415 0 0 $X=111425 $Y=112665
X429 1 2 9 dpp20_CDNS_724655180287 $T=163730 200845 0 90 $X=102650 $Y=189765
X430 1 2 9 dpp20_CDNS_724655180287 $T=241095 201100 0 90 $X=180015 $Y=190020
X431 2 3 1 rpp1k1_3_CDNS_724655180288 $T=16595 197030 0 0 $X=13435 $Y=196810
X432 15 14 1 rpp1k1_3_CDNS_724655180288 $T=56660 175685 0 0 $X=53500 $Y=175465
X433 5 6 11 1 pe3_CDNS_724655180289 $T=20540 115965 1 0 $X=19030 $Y=114495
X434 5 7 12 1 pe3_CDNS_724655180289 $T=23860 115965 1 0 $X=22350 $Y=114495
X435 5 12 13 1 pe3_CDNS_724655180289 $T=27180 115965 1 0 $X=25670 $Y=114495
X436 2 MASCO__X4 $T=376810 225310 0 0 $X=376810 $Y=225310
X437 2 MASCO__X4 $T=378810 225310 0 0 $X=378810 $Y=225310
X438 2 MASCO__X4 $T=380810 225310 0 0 $X=380810 $Y=225310
X439 2 MASCO__X4 $T=382810 225310 0 0 $X=382810 $Y=225310
X440 2 MASCO__X4 $T=384810 225310 0 0 $X=384810 $Y=225310
X441 9 MASCO__X4 $T=385495 160110 0 0 $X=385495 $Y=160110
X442 2 MASCO__X4 $T=386810 225310 0 0 $X=386810 $Y=225310
X443 9 MASCO__X4 $T=387495 160110 0 0 $X=387495 $Y=160110
X444 2 MASCO__X4 $T=388810 225310 0 0 $X=388810 $Y=225310
X445 9 MASCO__X4 $T=389495 160110 0 0 $X=389495 $Y=160110
X446 2 MASCO__X4 $T=390810 225310 0 0 $X=390810 $Y=225310
X447 9 MASCO__X4 $T=391495 160110 0 0 $X=391495 $Y=160110
X448 2 MASCO__X4 $T=392810 225310 0 0 $X=392810 $Y=225310
X449 9 MASCO__X4 $T=393495 160110 0 0 $X=393495 $Y=160110
X450 2 MASCO__X4 $T=394810 225310 0 0 $X=394810 $Y=225310
X451 9 MASCO__X4 $T=395495 160110 0 0 $X=395495 $Y=160110
X452 2 MASCO__X4 $T=396810 225310 0 0 $X=396810 $Y=225310
X453 9 MASCO__X4 $T=397495 160110 0 0 $X=397495 $Y=160110
X454 2 MASCO__X4 $T=398810 225310 0 0 $X=398810 $Y=225310
X455 9 MASCO__X4 $T=399495 160110 0 0 $X=399495 $Y=160110
X456 2 MASCO__X4 $T=400810 225310 0 0 $X=400810 $Y=225310
X457 9 MASCO__X4 $T=401495 160110 0 0 $X=401495 $Y=160110
X458 2 MASCO__X4 $T=402810 225310 0 0 $X=402810 $Y=225310
X459 9 MASCO__X4 $T=403495 160110 0 0 $X=403495 $Y=160110
X460 2 MASCO__X5 $T=376810 211310 0 0 $X=376810 $Y=211310
X461 2 MASCO__X5 $T=378810 211310 0 0 $X=378810 $Y=211310
X462 2 MASCO__X5 $T=380810 211310 0 0 $X=380810 $Y=211310
X463 2 MASCO__X5 $T=382810 211310 0 0 $X=382810 $Y=211310
X464 2 MASCO__X5 $T=384810 211310 0 0 $X=384810 $Y=211310
X465 9 MASCO__X5 $T=385495 146110 0 0 $X=385495 $Y=146110
X466 2 MASCO__X5 $T=386810 211310 0 0 $X=386810 $Y=211310
X467 9 MASCO__X5 $T=387495 146110 0 0 $X=387495 $Y=146110
X468 2 MASCO__X5 $T=388810 211310 0 0 $X=388810 $Y=211310
X469 9 MASCO__X5 $T=389495 146110 0 0 $X=389495 $Y=146110
X470 2 MASCO__X5 $T=390810 211310 0 0 $X=390810 $Y=211310
X471 9 MASCO__X5 $T=391495 146110 0 0 $X=391495 $Y=146110
X472 2 MASCO__X5 $T=392810 211310 0 0 $X=392810 $Y=211310
X473 9 MASCO__X5 $T=393495 146110 0 0 $X=393495 $Y=146110
X474 2 MASCO__X5 $T=394810 211310 0 0 $X=394810 $Y=211310
X475 9 MASCO__X5 $T=395495 146110 0 0 $X=395495 $Y=146110
X476 2 MASCO__X5 $T=396810 211310 0 0 $X=396810 $Y=211310
X477 9 MASCO__X5 $T=397495 146110 0 0 $X=397495 $Y=146110
X478 2 MASCO__X5 $T=398810 211310 0 0 $X=398810 $Y=211310
X479 9 MASCO__X5 $T=399495 146110 0 0 $X=399495 $Y=146110
X480 2 MASCO__X5 $T=400810 211310 0 0 $X=400810 $Y=211310
X481 9 MASCO__X5 $T=401495 146110 0 0 $X=401495 $Y=146110
X482 2 MASCO__X5 $T=402810 211310 0 0 $X=402810 $Y=211310
X483 9 MASCO__X5 $T=403495 146110 0 0 $X=403495 $Y=146110
X484 9 MASCO__X6 $T=234495 155110 0 0 $X=234495 $Y=155110
X485 9 MASCO__X6 $T=236495 155110 0 0 $X=236495 $Y=155110
X486 9 MASCO__X6 $T=238495 155110 0 0 $X=238495 $Y=155110
X487 9 MASCO__X6 $T=240495 155110 0 0 $X=240495 $Y=155110
X488 9 MASCO__X6 $T=242495 155110 0 0 $X=242495 $Y=155110
X489 9 MASCO__X6 $T=244495 155110 0 0 $X=244495 $Y=155110
X490 9 MASCO__X6 $T=246495 155110 0 0 $X=246495 $Y=155110
X491 9 MASCO__X6 $T=248495 155110 0 0 $X=248495 $Y=155110
X492 9 MASCO__X6 $T=250495 155110 0 0 $X=250495 $Y=155110
X493 9 MASCO__X6 $T=252495 155110 0 0 $X=252495 $Y=155110
X494 9 MASCO__X6 $T=254495 155110 0 0 $X=254495 $Y=155110
X495 9 MASCO__X6 $T=256495 155110 0 0 $X=256495 $Y=155110
X496 9 MASCO__X6 $T=258495 155110 0 0 $X=258495 $Y=155110
X497 9 MASCO__X6 $T=260495 155110 0 0 $X=260495 $Y=155110
X498 9 MASCO__X6 $T=262495 155110 0 0 $X=262495 $Y=155110
X499 9 MASCO__X6 $T=264495 155110 0 0 $X=264495 $Y=155110
X500 9 MASCO__X6 $T=266495 155110 0 0 $X=266495 $Y=155110
X501 9 MASCO__X6 $T=270495 155110 0 0 $X=270495 $Y=155110
X502 9 MASCO__X6 $T=272495 155110 0 0 $X=272495 $Y=155110
X503 9 MASCO__X6 $T=274495 155110 0 0 $X=274495 $Y=155110
X504 9 MASCO__X6 $T=276495 155110 0 0 $X=276495 $Y=155110
X505 9 MASCO__X6 $T=278495 155110 0 0 $X=278495 $Y=155110
X506 9 MASCO__X6 $T=280495 155110 0 0 $X=280495 $Y=155110
X507 9 MASCO__X6 $T=282495 155110 0 0 $X=282495 $Y=155110
X508 9 MASCO__X6 $T=284495 155110 0 0 $X=284495 $Y=155110
X509 9 MASCO__X6 $T=286495 155110 0 0 $X=286495 $Y=155110
X510 9 MASCO__X6 $T=288495 155110 0 0 $X=288495 $Y=155110
X511 9 MASCO__X6 $T=290495 155110 0 0 $X=290495 $Y=155110
X512 9 MASCO__X6 $T=292495 155110 0 0 $X=292495 $Y=155110
X513 9 MASCO__X6 $T=294495 155110 0 0 $X=294495 $Y=155110
X514 9 MASCO__X6 $T=296495 155110 0 0 $X=296495 $Y=155110
X515 9 MASCO__X6 $T=298495 155110 0 0 $X=298495 $Y=155110
X516 9 MASCO__X6 $T=300495 155110 0 0 $X=300495 $Y=155110
X517 9 MASCO__X6 $T=302495 155110 0 0 $X=302495 $Y=155110
X518 9 MASCO__X6 $T=304495 155110 0 0 $X=304495 $Y=155110
X519 9 MASCO__X6 $T=306495 155110 0 0 $X=306495 $Y=155110
X520 9 MASCO__X6 $T=308495 155110 0 0 $X=308495 $Y=155110
X521 9 MASCO__X6 $T=310495 155110 0 0 $X=310495 $Y=155110
X522 9 MASCO__X6 $T=312495 155110 0 0 $X=312495 $Y=155110
X523 9 MASCO__X6 $T=314495 155110 0 0 $X=314495 $Y=155110
X524 9 MASCO__X6 $T=316495 155110 0 0 $X=316495 $Y=155110
X525 9 MASCO__X6 $T=318495 155110 0 0 $X=318495 $Y=155110
X526 9 MASCO__X6 $T=320495 155110 0 0 $X=320495 $Y=155110
X527 9 MASCO__X6 $T=322495 155110 0 0 $X=322495 $Y=155110
X528 9 MASCO__X6 $T=324495 155110 0 0 $X=324495 $Y=155110
X529 9 MASCO__X6 $T=326495 155110 0 0 $X=326495 $Y=155110
X530 9 MASCO__X6 $T=328495 155110 0 0 $X=328495 $Y=155110
X531 9 MASCO__X6 $T=330495 155110 0 0 $X=330495 $Y=155110
X532 9 MASCO__X6 $T=332495 155110 0 0 $X=332495 $Y=155110
X533 9 MASCO__X6 $T=334495 155110 0 0 $X=334495 $Y=155110
X534 9 MASCO__X6 $T=336495 155110 0 0 $X=336495 $Y=155110
X535 9 MASCO__X6 $T=338495 155110 0 0 $X=338495 $Y=155110
X536 9 MASCO__X6 $T=340495 155110 0 0 $X=340495 $Y=155110
X537 9 MASCO__X6 $T=342495 155110 0 0 $X=342495 $Y=155110
X538 9 MASCO__X6 $T=344495 155110 0 0 $X=344495 $Y=155110
X539 9 MASCO__X6 $T=346495 155110 0 0 $X=346495 $Y=155110
X540 9 MASCO__X6 $T=348495 155110 0 0 $X=348495 $Y=155110
X541 9 MASCO__X6 $T=350495 155110 0 0 $X=350495 $Y=155110
X542 9 MASCO__X6 $T=352495 155110 0 0 $X=352495 $Y=155110
X543 9 MASCO__X6 $T=354495 155110 0 0 $X=354495 $Y=155110
X544 9 MASCO__X6 $T=356495 155110 0 0 $X=356495 $Y=155110
X545 9 MASCO__X6 $T=358495 155110 0 0 $X=358495 $Y=155110
X546 9 MASCO__X6 $T=360495 155110 0 0 $X=360495 $Y=155110
X547 9 MASCO__X6 $T=362495 155110 0 0 $X=362495 $Y=155110
X548 9 MASCO__X6 $T=364495 155110 0 0 $X=364495 $Y=155110
X549 9 MASCO__X6 $T=366495 155110 0 0 $X=366495 $Y=155110
X550 9 MASCO__X6 $T=368495 155110 0 0 $X=368495 $Y=155110
X551 9 MASCO__X6 $T=370495 155110 0 0 $X=370495 $Y=155110
X552 9 MASCO__X6 $T=372495 155110 0 0 $X=372495 $Y=155110
X553 2 MASCO__X6 $T=373810 210310 0 0 $X=373810 $Y=210310
X554 2 MASCO__X6 $T=373810 219310 0 0 $X=373810 $Y=219310
X555 9 MASCO__X6 $T=374495 155110 0 0 $X=374495 $Y=155110
X556 2 MASCO__X6 $T=377810 210310 0 0 $X=377810 $Y=210310
X557 2 MASCO__X6 $T=377810 219310 0 0 $X=377810 $Y=219310
X558 2 MASCO__X6 $T=377810 228310 0 0 $X=377810 $Y=228310
X559 2 MASCO__X6 $T=379810 210310 0 0 $X=379810 $Y=210310
X560 2 MASCO__X6 $T=379810 219310 0 0 $X=379810 $Y=219310
X561 2 MASCO__X6 $T=379810 228310 0 0 $X=379810 $Y=228310
X562 2 MASCO__X6 $T=381810 210310 0 0 $X=381810 $Y=210310
X563 2 MASCO__X6 $T=381810 219310 0 0 $X=381810 $Y=219310
X564 2 MASCO__X6 $T=381810 228310 0 0 $X=381810 $Y=228310
X565 2 MASCO__X6 $T=383810 210310 0 0 $X=383810 $Y=210310
X566 2 MASCO__X6 $T=383810 219310 0 0 $X=383810 $Y=219310
X567 2 MASCO__X6 $T=383810 228310 0 0 $X=383810 $Y=228310
X568 2 MASCO__X6 $T=385810 210310 0 0 $X=385810 $Y=210310
X569 2 MASCO__X6 $T=385810 219310 0 0 $X=385810 $Y=219310
X570 2 MASCO__X6 $T=385810 228310 0 0 $X=385810 $Y=228310
X571 9 MASCO__X6 $T=386495 145110 0 0 $X=386495 $Y=145110
X572 9 MASCO__X6 $T=386495 154110 0 0 $X=386495 $Y=154110
X573 9 MASCO__X6 $T=386495 163110 0 0 $X=386495 $Y=163110
X574 2 MASCO__X6 $T=387810 210310 0 0 $X=387810 $Y=210310
X575 2 MASCO__X6 $T=387810 219310 0 0 $X=387810 $Y=219310
X576 2 MASCO__X6 $T=387810 228310 0 0 $X=387810 $Y=228310
X577 9 MASCO__X6 $T=388495 145110 0 0 $X=388495 $Y=145110
X578 9 MASCO__X6 $T=388495 154110 0 0 $X=388495 $Y=154110
X579 9 MASCO__X6 $T=388495 163110 0 0 $X=388495 $Y=163110
X580 2 MASCO__X6 $T=389810 210310 0 0 $X=389810 $Y=210310
X581 2 MASCO__X6 $T=389810 219310 0 0 $X=389810 $Y=219310
X582 2 MASCO__X6 $T=389810 228310 0 0 $X=389810 $Y=228310
X583 9 MASCO__X6 $T=390495 145110 0 0 $X=390495 $Y=145110
X584 9 MASCO__X6 $T=390495 154110 0 0 $X=390495 $Y=154110
X585 9 MASCO__X6 $T=390495 163110 0 0 $X=390495 $Y=163110
X586 2 MASCO__X6 $T=391810 210310 0 0 $X=391810 $Y=210310
X587 2 MASCO__X6 $T=391810 219310 0 0 $X=391810 $Y=219310
X588 2 MASCO__X6 $T=391810 228310 0 0 $X=391810 $Y=228310
X589 9 MASCO__X6 $T=392495 145110 0 0 $X=392495 $Y=145110
X590 9 MASCO__X6 $T=392495 154110 0 0 $X=392495 $Y=154110
X591 9 MASCO__X6 $T=392495 163110 0 0 $X=392495 $Y=163110
X592 2 MASCO__X6 $T=393810 210310 0 0 $X=393810 $Y=210310
X593 2 MASCO__X6 $T=393810 219310 0 0 $X=393810 $Y=219310
X594 2 MASCO__X6 $T=393810 228310 0 0 $X=393810 $Y=228310
X595 9 MASCO__X6 $T=394495 145110 0 0 $X=394495 $Y=145110
X596 9 MASCO__X6 $T=394495 154110 0 0 $X=394495 $Y=154110
X597 9 MASCO__X6 $T=394495 163110 0 0 $X=394495 $Y=163110
X598 2 MASCO__X6 $T=395810 210310 0 0 $X=395810 $Y=210310
X599 2 MASCO__X6 $T=395810 219310 0 0 $X=395810 $Y=219310
X600 2 MASCO__X6 $T=395810 228310 0 0 $X=395810 $Y=228310
X601 9 MASCO__X6 $T=396495 145110 0 0 $X=396495 $Y=145110
X602 9 MASCO__X6 $T=396495 154110 0 0 $X=396495 $Y=154110
X603 9 MASCO__X6 $T=396495 163110 0 0 $X=396495 $Y=163110
X604 2 MASCO__X6 $T=397810 210310 0 0 $X=397810 $Y=210310
X605 2 MASCO__X6 $T=397810 219310 0 0 $X=397810 $Y=219310
X606 2 MASCO__X6 $T=397810 228310 0 0 $X=397810 $Y=228310
X607 9 MASCO__X6 $T=398495 145110 0 0 $X=398495 $Y=145110
X608 9 MASCO__X6 $T=398495 154110 0 0 $X=398495 $Y=154110
X609 9 MASCO__X6 $T=398495 163110 0 0 $X=398495 $Y=163110
X610 2 MASCO__X6 $T=399810 210310 0 0 $X=399810 $Y=210310
X611 2 MASCO__X6 $T=399810 219310 0 0 $X=399810 $Y=219310
X612 2 MASCO__X6 $T=399810 228310 0 0 $X=399810 $Y=228310
X613 9 MASCO__X6 $T=400495 145110 0 0 $X=400495 $Y=145110
X614 9 MASCO__X6 $T=400495 154110 0 0 $X=400495 $Y=154110
X615 9 MASCO__X6 $T=400495 163110 0 0 $X=400495 $Y=163110
X616 2 MASCO__X6 $T=401810 210310 0 0 $X=401810 $Y=210310
X617 2 MASCO__X6 $T=401810 219310 0 0 $X=401810 $Y=219310
X618 2 MASCO__X6 $T=401810 228310 0 0 $X=401810 $Y=228310
X619 9 MASCO__X6 $T=402495 145110 0 0 $X=402495 $Y=145110
X620 9 MASCO__X6 $T=402495 154110 0 0 $X=402495 $Y=154110
X621 9 MASCO__X6 $T=402495 163110 0 0 $X=402495 $Y=163110
X622 9 MASCO__X7 $T=234495 164110 0 0 $X=234495 $Y=164110
X623 9 MASCO__X7 $T=236495 164110 0 0 $X=236495 $Y=164110
X624 9 MASCO__X7 $T=238495 164110 0 0 $X=238495 $Y=164110
X625 9 MASCO__X7 $T=240495 164110 0 0 $X=240495 $Y=164110
X626 9 MASCO__X7 $T=242495 164110 0 0 $X=242495 $Y=164110
X627 9 MASCO__X7 $T=244495 164110 0 0 $X=244495 $Y=164110
X628 9 MASCO__X7 $T=246495 164110 0 0 $X=246495 $Y=164110
X629 9 MASCO__X7 $T=248495 164110 0 0 $X=248495 $Y=164110
X630 9 MASCO__X7 $T=250495 164110 0 0 $X=250495 $Y=164110
X631 9 MASCO__X7 $T=252495 164110 0 0 $X=252495 $Y=164110
X632 9 MASCO__X7 $T=254495 164110 0 0 $X=254495 $Y=164110
X633 9 MASCO__X7 $T=256495 164110 0 0 $X=256495 $Y=164110
X634 9 MASCO__X7 $T=258495 164110 0 0 $X=258495 $Y=164110
X635 9 MASCO__X7 $T=260495 164110 0 0 $X=260495 $Y=164110
X636 9 MASCO__X7 $T=262495 164110 0 0 $X=262495 $Y=164110
X637 9 MASCO__X7 $T=264495 164110 0 0 $X=264495 $Y=164110
X638 9 MASCO__X7 $T=266495 164110 0 0 $X=266495 $Y=164110
X639 9 MASCO__X7 $T=270495 164110 0 0 $X=270495 $Y=164110
X640 9 MASCO__X7 $T=272495 164110 0 0 $X=272495 $Y=164110
X641 9 MASCO__X7 $T=274495 164110 0 0 $X=274495 $Y=164110
X642 9 MASCO__X7 $T=276495 164110 0 0 $X=276495 $Y=164110
X643 9 MASCO__X7 $T=278495 164110 0 0 $X=278495 $Y=164110
X644 9 MASCO__X7 $T=280495 164110 0 0 $X=280495 $Y=164110
X645 9 MASCO__X7 $T=282495 164110 0 0 $X=282495 $Y=164110
X646 9 MASCO__X7 $T=284495 164110 0 0 $X=284495 $Y=164110
X647 9 MASCO__X7 $T=286495 164110 0 0 $X=286495 $Y=164110
X648 9 MASCO__X7 $T=288495 164110 0 0 $X=288495 $Y=164110
X649 9 MASCO__X7 $T=290495 164110 0 0 $X=290495 $Y=164110
X650 9 MASCO__X7 $T=292495 164110 0 0 $X=292495 $Y=164110
X651 9 MASCO__X7 $T=294495 164110 0 0 $X=294495 $Y=164110
X652 9 MASCO__X7 $T=296495 164110 0 0 $X=296495 $Y=164110
X653 9 MASCO__X7 $T=298495 164110 0 0 $X=298495 $Y=164110
X654 9 MASCO__X7 $T=300495 164110 0 0 $X=300495 $Y=164110
X655 9 MASCO__X7 $T=302495 164110 0 0 $X=302495 $Y=164110
X656 9 MASCO__X7 $T=304495 164110 0 0 $X=304495 $Y=164110
X657 9 MASCO__X7 $T=306495 164110 0 0 $X=306495 $Y=164110
X658 9 MASCO__X7 $T=308495 164110 0 0 $X=308495 $Y=164110
X659 9 MASCO__X7 $T=310495 164110 0 0 $X=310495 $Y=164110
X660 9 MASCO__X7 $T=312495 164110 0 0 $X=312495 $Y=164110
X661 9 MASCO__X7 $T=314495 164110 0 0 $X=314495 $Y=164110
X662 9 MASCO__X7 $T=316495 164110 0 0 $X=316495 $Y=164110
X663 9 MASCO__X7 $T=318495 164110 0 0 $X=318495 $Y=164110
X664 9 MASCO__X7 $T=320495 164110 0 0 $X=320495 $Y=164110
X665 9 MASCO__X7 $T=322495 164110 0 0 $X=322495 $Y=164110
X666 9 MASCO__X7 $T=324495 164110 0 0 $X=324495 $Y=164110
X667 9 MASCO__X7 $T=326495 164110 0 0 $X=326495 $Y=164110
X668 9 MASCO__X7 $T=328495 164110 0 0 $X=328495 $Y=164110
X669 9 MASCO__X7 $T=330495 164110 0 0 $X=330495 $Y=164110
X670 9 MASCO__X7 $T=332495 164110 0 0 $X=332495 $Y=164110
X671 9 MASCO__X7 $T=334495 164110 0 0 $X=334495 $Y=164110
X672 9 MASCO__X7 $T=336495 164110 0 0 $X=336495 $Y=164110
X673 9 MASCO__X7 $T=338495 164110 0 0 $X=338495 $Y=164110
X674 9 MASCO__X7 $T=340495 164110 0 0 $X=340495 $Y=164110
X675 9 MASCO__X7 $T=342495 164110 0 0 $X=342495 $Y=164110
X676 9 MASCO__X7 $T=344495 164110 0 0 $X=344495 $Y=164110
X677 9 MASCO__X7 $T=346495 164110 0 0 $X=346495 $Y=164110
X678 9 MASCO__X7 $T=348495 164110 0 0 $X=348495 $Y=164110
X679 9 MASCO__X7 $T=350495 164110 0 0 $X=350495 $Y=164110
X680 9 MASCO__X7 $T=352495 164110 0 0 $X=352495 $Y=164110
X681 9 MASCO__X7 $T=354495 164110 0 0 $X=354495 $Y=164110
X682 9 MASCO__X7 $T=356495 164110 0 0 $X=356495 $Y=164110
X683 9 MASCO__X7 $T=358495 164110 0 0 $X=358495 $Y=164110
X684 9 MASCO__X7 $T=360495 164110 0 0 $X=360495 $Y=164110
X685 9 MASCO__X7 $T=362495 164110 0 0 $X=362495 $Y=164110
X686 9 MASCO__X7 $T=364495 164110 0 0 $X=364495 $Y=164110
X687 9 MASCO__X7 $T=366495 164110 0 0 $X=366495 $Y=164110
X688 9 MASCO__X7 $T=368495 164110 0 0 $X=368495 $Y=164110
X689 9 MASCO__X7 $T=370495 164110 0 0 $X=370495 $Y=164110
X690 9 MASCO__X7 $T=372495 164110 0 0 $X=372495 $Y=164110
X691 9 MASCO__X7 $T=374495 164110 0 0 $X=374495 $Y=164110
X692 9 MASCO__X7 $T=378495 164110 0 0 $X=378495 $Y=164110
X693 9 MASCO__X7 $T=380495 164110 0 0 $X=380495 $Y=164110
X694 9 MASCO__X7 $T=382495 164110 0 0 $X=382495 $Y=164110
X695 9 MASCO__X7 $T=384495 164110 0 0 $X=384495 $Y=164110
X696 9 MASCO__X8 $T=233495 156110 0 0 $X=233495 $Y=156110
X697 9 MASCO__X8 $T=235495 156110 0 0 $X=235495 $Y=156110
X698 9 MASCO__X8 $T=237495 156110 0 0 $X=237495 $Y=156110
X699 9 MASCO__X8 $T=239495 156110 0 0 $X=239495 $Y=156110
X700 9 MASCO__X8 $T=241495 156110 0 0 $X=241495 $Y=156110
X701 9 MASCO__X8 $T=243495 156110 0 0 $X=243495 $Y=156110
X702 9 MASCO__X8 $T=245495 156110 0 0 $X=245495 $Y=156110
X703 9 MASCO__X8 $T=247495 156110 0 0 $X=247495 $Y=156110
X704 9 MASCO__X8 $T=249495 156110 0 0 $X=249495 $Y=156110
X705 9 MASCO__X8 $T=251495 156110 0 0 $X=251495 $Y=156110
X706 9 MASCO__X8 $T=253495 156110 0 0 $X=253495 $Y=156110
X707 9 MASCO__X8 $T=255495 156110 0 0 $X=255495 $Y=156110
X708 9 MASCO__X8 $T=257495 156110 0 0 $X=257495 $Y=156110
X709 9 MASCO__X8 $T=259495 156110 0 0 $X=259495 $Y=156110
X710 9 MASCO__X8 $T=261495 156110 0 0 $X=261495 $Y=156110
X711 9 MASCO__X8 $T=263495 156110 0 0 $X=263495 $Y=156110
X712 9 MASCO__X8 $T=265495 156110 0 0 $X=265495 $Y=156110
X713 9 MASCO__X8 $T=269495 156110 0 0 $X=269495 $Y=156110
X714 9 MASCO__X8 $T=271495 156110 0 0 $X=271495 $Y=156110
X715 9 MASCO__X8 $T=273495 156110 0 0 $X=273495 $Y=156110
X716 9 MASCO__X8 $T=275495 156110 0 0 $X=275495 $Y=156110
X717 9 MASCO__X8 $T=277495 156110 0 0 $X=277495 $Y=156110
X718 9 MASCO__X8 $T=279495 156110 0 0 $X=279495 $Y=156110
X719 9 MASCO__X8 $T=281495 156110 0 0 $X=281495 $Y=156110
X720 9 MASCO__X8 $T=283495 156110 0 0 $X=283495 $Y=156110
X721 9 MASCO__X8 $T=285495 156110 0 0 $X=285495 $Y=156110
X722 9 MASCO__X8 $T=287495 156110 0 0 $X=287495 $Y=156110
X723 9 MASCO__X8 $T=289495 156110 0 0 $X=289495 $Y=156110
X724 9 MASCO__X8 $T=291495 156110 0 0 $X=291495 $Y=156110
X725 9 MASCO__X8 $T=293495 156110 0 0 $X=293495 $Y=156110
X726 9 MASCO__X8 $T=295495 156110 0 0 $X=295495 $Y=156110
X727 9 MASCO__X8 $T=297495 156110 0 0 $X=297495 $Y=156110
X728 9 MASCO__X8 $T=299495 156110 0 0 $X=299495 $Y=156110
X729 9 MASCO__X8 $T=301495 156110 0 0 $X=301495 $Y=156110
X730 9 MASCO__X8 $T=303495 156110 0 0 $X=303495 $Y=156110
X731 9 MASCO__X8 $T=305495 156110 0 0 $X=305495 $Y=156110
X732 9 MASCO__X8 $T=307495 156110 0 0 $X=307495 $Y=156110
X733 9 MASCO__X8 $T=309495 156110 0 0 $X=309495 $Y=156110
X734 9 MASCO__X8 $T=311495 156110 0 0 $X=311495 $Y=156110
X735 9 MASCO__X8 $T=313495 156110 0 0 $X=313495 $Y=156110
X736 9 MASCO__X8 $T=315495 156110 0 0 $X=315495 $Y=156110
X737 9 MASCO__X8 $T=317495 156110 0 0 $X=317495 $Y=156110
X738 9 MASCO__X8 $T=319495 156110 0 0 $X=319495 $Y=156110
X739 9 MASCO__X8 $T=321495 156110 0 0 $X=321495 $Y=156110
X740 9 MASCO__X8 $T=323495 156110 0 0 $X=323495 $Y=156110
X741 9 MASCO__X8 $T=325495 156110 0 0 $X=325495 $Y=156110
X742 9 MASCO__X8 $T=327495 156110 0 0 $X=327495 $Y=156110
X743 9 MASCO__X8 $T=329495 156110 0 0 $X=329495 $Y=156110
X744 9 MASCO__X8 $T=331495 156110 0 0 $X=331495 $Y=156110
X745 9 MASCO__X8 $T=333495 156110 0 0 $X=333495 $Y=156110
X746 9 MASCO__X8 $T=335495 156110 0 0 $X=335495 $Y=156110
X747 9 MASCO__X8 $T=337495 156110 0 0 $X=337495 $Y=156110
X748 9 MASCO__X8 $T=339495 156110 0 0 $X=339495 $Y=156110
X749 9 MASCO__X8 $T=341495 156110 0 0 $X=341495 $Y=156110
X750 9 MASCO__X8 $T=343495 156110 0 0 $X=343495 $Y=156110
X751 9 MASCO__X8 $T=345495 156110 0 0 $X=345495 $Y=156110
X752 9 MASCO__X8 $T=347495 156110 0 0 $X=347495 $Y=156110
X753 9 MASCO__X8 $T=349495 156110 0 0 $X=349495 $Y=156110
X754 9 MASCO__X8 $T=351495 156110 0 0 $X=351495 $Y=156110
X755 9 MASCO__X8 $T=353495 156110 0 0 $X=353495 $Y=156110
X756 9 MASCO__X8 $T=355495 156110 0 0 $X=355495 $Y=156110
X757 9 MASCO__X8 $T=357495 156110 0 0 $X=357495 $Y=156110
X758 9 MASCO__X8 $T=359495 156110 0 0 $X=359495 $Y=156110
X759 9 MASCO__X8 $T=361495 156110 0 0 $X=361495 $Y=156110
X760 9 MASCO__X8 $T=363495 156110 0 0 $X=363495 $Y=156110
X761 9 MASCO__X8 $T=365495 156110 0 0 $X=365495 $Y=156110
X762 9 MASCO__X8 $T=367495 156110 0 0 $X=367495 $Y=156110
X763 9 MASCO__X8 $T=369495 156110 0 0 $X=369495 $Y=156110
X764 9 MASCO__X8 $T=371495 156110 0 0 $X=371495 $Y=156110
X765 9 MASCO__X8 $T=373495 156110 0 0 $X=373495 $Y=156110
X766 9 MASCO__X8 $T=377495 156110 0 0 $X=377495 $Y=156110
X767 9 MASCO__X8 $T=379495 156110 0 0 $X=379495 $Y=156110
X768 9 MASCO__X8 $T=381495 156110 0 0 $X=381495 $Y=156110
X769 9 MASCO__X8 $T=383495 156110 0 0 $X=383495 $Y=156110
X770 2 MASCO__X10 $T=271810 218310 0 0 $X=271810 $Y=218310
X771 2 MASCO__X10 $T=273810 218310 0 0 $X=273810 $Y=218310
X772 2 MASCO__X10 $T=275810 218310 0 0 $X=275810 $Y=218310
X773 2 MASCO__X10 $T=277810 218310 0 0 $X=277810 $Y=218310
X774 2 MASCO__X10 $T=279810 218310 0 0 $X=279810 $Y=218310
X775 2 MASCO__X10 $T=281810 218310 0 0 $X=281810 $Y=218310
X776 2 MASCO__X10 $T=283810 218310 0 0 $X=283810 $Y=218310
X777 2 MASCO__X10 $T=285810 218310 0 0 $X=285810 $Y=218310
X778 2 MASCO__X10 $T=287810 218310 0 0 $X=287810 $Y=218310
X779 2 MASCO__X10 $T=289810 218310 0 0 $X=289810 $Y=218310
X780 2 MASCO__X10 $T=291810 218310 0 0 $X=291810 $Y=218310
X781 2 MASCO__X10 $T=293810 218310 0 0 $X=293810 $Y=218310
X782 2 MASCO__X10 $T=295810 218310 0 0 $X=295810 $Y=218310
X783 2 MASCO__X10 $T=297810 218310 0 0 $X=297810 $Y=218310
X784 2 MASCO__X10 $T=299810 218310 0 0 $X=299810 $Y=218310
X785 2 MASCO__X10 $T=301810 218310 0 0 $X=301810 $Y=218310
X786 2 MASCO__X10 $T=303810 218310 0 0 $X=303810 $Y=218310
X787 2 MASCO__X10 $T=305810 218310 0 0 $X=305810 $Y=218310
X788 2 MASCO__X10 $T=307810 218310 0 0 $X=307810 $Y=218310
X789 2 MASCO__X10 $T=309810 218310 0 0 $X=309810 $Y=218310
X790 2 MASCO__X10 $T=311810 218310 0 0 $X=311810 $Y=218310
X791 2 MASCO__X10 $T=313810 218310 0 0 $X=313810 $Y=218310
X792 2 MASCO__X10 $T=315810 218310 0 0 $X=315810 $Y=218310
X793 2 MASCO__X10 $T=317810 218310 0 0 $X=317810 $Y=218310
X794 2 MASCO__X10 $T=319810 218310 0 0 $X=319810 $Y=218310
X795 2 MASCO__X10 $T=321810 218310 0 0 $X=321810 $Y=218310
X796 2 MASCO__X10 $T=323810 218310 0 0 $X=323810 $Y=218310
X797 2 MASCO__X10 $T=325810 218310 0 0 $X=325810 $Y=218310
X798 2 MASCO__X10 $T=327810 218310 0 0 $X=327810 $Y=218310
X799 2 MASCO__X10 $T=329810 218310 0 0 $X=329810 $Y=218310
X800 2 MASCO__X10 $T=331810 218310 0 0 $X=331810 $Y=218310
X801 2 MASCO__X10 $T=333810 218310 0 0 $X=333810 $Y=218310
X802 2 MASCO__X10 $T=335810 218310 0 0 $X=335810 $Y=218310
X803 2 MASCO__X10 $T=337810 218310 0 0 $X=337810 $Y=218310
X804 2 MASCO__X10 $T=339810 218310 0 0 $X=339810 $Y=218310
X805 2 MASCO__X10 $T=341810 218310 0 0 $X=341810 $Y=218310
X806 2 MASCO__X10 $T=343810 218310 0 0 $X=343810 $Y=218310
X807 2 MASCO__X10 $T=345810 218310 0 0 $X=345810 $Y=218310
X808 2 MASCO__X10 $T=347810 218310 0 0 $X=347810 $Y=218310
X809 2 MASCO__X10 $T=349810 218310 0 0 $X=349810 $Y=218310
X810 2 MASCO__X10 $T=351810 218310 0 0 $X=351810 $Y=218310
X811 2 MASCO__X10 $T=353810 218310 0 0 $X=353810 $Y=218310
X812 2 MASCO__X10 $T=355810 218310 0 0 $X=355810 $Y=218310
X813 2 MASCO__X10 $T=357810 218310 0 0 $X=357810 $Y=218310
X814 2 MASCO__X10 $T=359810 218310 0 0 $X=359810 $Y=218310
X815 2 MASCO__X10 $T=361810 218310 0 0 $X=361810 $Y=218310
X816 2 MASCO__X10 $T=363810 218310 0 0 $X=363810 $Y=218310
X817 2 MASCO__X10 $T=365810 218310 0 0 $X=365810 $Y=218310
X818 2 MASCO__X10 $T=367810 218310 0 0 $X=367810 $Y=218310
X819 2 MASCO__X10 $T=369810 218310 0 0 $X=369810 $Y=218310
X820 2 MASCO__X10 $T=371810 218310 0 0 $X=371810 $Y=218310
X821 2 MASCO__X11 $T=271810 210310 0 0 $X=271810 $Y=210310
X822 2 MASCO__X11 $T=273810 210310 0 0 $X=273810 $Y=210310
X823 2 MASCO__X11 $T=275810 210310 0 0 $X=275810 $Y=210310
X824 2 MASCO__X11 $T=277810 210310 0 0 $X=277810 $Y=210310
X825 2 MASCO__X11 $T=279810 210310 0 0 $X=279810 $Y=210310
X826 2 MASCO__X11 $T=281810 210310 0 0 $X=281810 $Y=210310
X827 2 MASCO__X11 $T=283810 210310 0 0 $X=283810 $Y=210310
X828 2 MASCO__X11 $T=285810 210310 0 0 $X=285810 $Y=210310
X829 2 MASCO__X11 $T=287810 210310 0 0 $X=287810 $Y=210310
X830 2 MASCO__X11 $T=289810 210310 0 0 $X=289810 $Y=210310
X831 2 MASCO__X11 $T=291810 210310 0 0 $X=291810 $Y=210310
X832 2 MASCO__X11 $T=293810 210310 0 0 $X=293810 $Y=210310
X833 2 MASCO__X11 $T=295810 210310 0 0 $X=295810 $Y=210310
X834 2 MASCO__X11 $T=297810 210310 0 0 $X=297810 $Y=210310
X835 2 MASCO__X11 $T=299810 210310 0 0 $X=299810 $Y=210310
X836 2 MASCO__X11 $T=301810 210310 0 0 $X=301810 $Y=210310
X837 2 MASCO__X11 $T=303810 210310 0 0 $X=303810 $Y=210310
X838 2 MASCO__X11 $T=305810 210310 0 0 $X=305810 $Y=210310
X839 2 MASCO__X11 $T=307810 210310 0 0 $X=307810 $Y=210310
X840 2 MASCO__X11 $T=309810 210310 0 0 $X=309810 $Y=210310
X841 2 MASCO__X11 $T=311810 210310 0 0 $X=311810 $Y=210310
X842 2 MASCO__X11 $T=313810 210310 0 0 $X=313810 $Y=210310
X843 2 MASCO__X11 $T=315810 210310 0 0 $X=315810 $Y=210310
X844 2 MASCO__X11 $T=317810 210310 0 0 $X=317810 $Y=210310
X845 2 MASCO__X11 $T=319810 210310 0 0 $X=319810 $Y=210310
X846 2 MASCO__X11 $T=321810 210310 0 0 $X=321810 $Y=210310
X847 2 MASCO__X11 $T=323810 210310 0 0 $X=323810 $Y=210310
X848 2 MASCO__X11 $T=325810 210310 0 0 $X=325810 $Y=210310
X849 2 MASCO__X11 $T=327810 210310 0 0 $X=327810 $Y=210310
X850 2 MASCO__X11 $T=329810 210310 0 0 $X=329810 $Y=210310
X851 2 MASCO__X11 $T=331810 210310 0 0 $X=331810 $Y=210310
X852 2 MASCO__X11 $T=333810 210310 0 0 $X=333810 $Y=210310
X853 2 MASCO__X11 $T=335810 210310 0 0 $X=335810 $Y=210310
X854 2 MASCO__X11 $T=337810 210310 0 0 $X=337810 $Y=210310
X855 2 MASCO__X11 $T=339810 210310 0 0 $X=339810 $Y=210310
X856 2 MASCO__X11 $T=341810 210310 0 0 $X=341810 $Y=210310
X857 2 MASCO__X11 $T=343810 210310 0 0 $X=343810 $Y=210310
X858 2 MASCO__X11 $T=345810 210310 0 0 $X=345810 $Y=210310
X859 2 MASCO__X11 $T=347810 210310 0 0 $X=347810 $Y=210310
X860 2 MASCO__X11 $T=349810 210310 0 0 $X=349810 $Y=210310
X861 2 MASCO__X11 $T=351810 210310 0 0 $X=351810 $Y=210310
X862 2 MASCO__X11 $T=353810 210310 0 0 $X=353810 $Y=210310
X863 2 MASCO__X11 $T=355810 210310 0 0 $X=355810 $Y=210310
X864 2 MASCO__X11 $T=357810 210310 0 0 $X=357810 $Y=210310
X865 2 MASCO__X11 $T=359810 210310 0 0 $X=359810 $Y=210310
X866 2 MASCO__X11 $T=361810 210310 0 0 $X=361810 $Y=210310
X867 2 MASCO__X11 $T=363810 210310 0 0 $X=363810 $Y=210310
X868 2 MASCO__X11 $T=365810 210310 0 0 $X=365810 $Y=210310
X869 2 MASCO__X11 $T=367810 210310 0 0 $X=367810 $Y=210310
X870 2 MASCO__X11 $T=369810 210310 0 0 $X=369810 $Y=210310
X871 2 MASCO__X11 $T=371810 210310 0 0 $X=371810 $Y=210310
X872 2 MASCO__Y13 $T=270810 219310 0 0 $X=270810 $Y=219310
X873 2 MASCO__Y13 $T=278810 219310 0 0 $X=278810 $Y=219310
X874 2 MASCO__Y13 $T=286810 219310 0 0 $X=286810 $Y=219310
X875 2 MASCO__Y13 $T=294810 219310 0 0 $X=294810 $Y=219310
X876 2 MASCO__Y13 $T=302810 219310 0 0 $X=302810 $Y=219310
X877 2 MASCO__Y13 $T=310810 219310 0 0 $X=310810 $Y=219310
X878 2 MASCO__Y13 $T=318810 219310 0 0 $X=318810 $Y=219310
X879 2 MASCO__Y13 $T=326810 219310 0 0 $X=326810 $Y=219310
X880 2 MASCO__Y13 $T=334810 219310 0 0 $X=334810 $Y=219310
X881 2 MASCO__Y13 $T=342810 219310 0 0 $X=342810 $Y=219310
X882 2 MASCO__Y13 $T=350810 219310 0 0 $X=350810 $Y=219310
X883 2 MASCO__Y13 $T=358810 219310 0 0 $X=358810 $Y=219310
X884 2 MASCO__Y13 $T=366810 219310 0 0 $X=366810 $Y=219310
X885 2 MASCO__Y14 $T=270810 237310 0 0 $X=270810 $Y=237310
X886 2 MASCO__Y14 $T=278810 237310 0 0 $X=278810 $Y=237310
X887 2 MASCO__Y14 $T=286810 237310 0 0 $X=286810 $Y=237310
X888 2 MASCO__Y14 $T=294810 237310 0 0 $X=294810 $Y=237310
X889 2 MASCO__Y14 $T=302810 237310 0 0 $X=302810 $Y=237310
X890 2 MASCO__Y14 $T=310810 237310 0 0 $X=310810 $Y=237310
X891 2 MASCO__Y14 $T=318810 237310 0 0 $X=318810 $Y=237310
X892 2 MASCO__Y14 $T=326810 237310 0 0 $X=326810 $Y=237310
X893 2 MASCO__Y14 $T=334810 237310 0 0 $X=334810 $Y=237310
X894 2 MASCO__Y14 $T=342810 237310 0 0 $X=342810 $Y=237310
X895 2 MASCO__Y14 $T=350810 237310 0 0 $X=350810 $Y=237310
X896 2 MASCO__Y14 $T=358810 237310 0 0 $X=358810 $Y=237310
X897 2 MASCO__Y14 $T=366810 237310 0 0 $X=366810 $Y=237310
X898 2 MASCO__Y15 $T=270810 211310 0 0 $X=270810 $Y=211310
X899 2 MASCO__Y15 $T=270810 213310 0 0 $X=270810 $Y=213310
X900 2 MASCO__Y15 $T=270810 215310 0 0 $X=270810 $Y=215310
X901 2 MASCO__Y15 $T=278810 211310 0 0 $X=278810 $Y=211310
X902 2 MASCO__Y15 $T=278810 213310 0 0 $X=278810 $Y=213310
X903 2 MASCO__Y15 $T=278810 215310 0 0 $X=278810 $Y=215310
X904 2 MASCO__Y15 $T=286810 211310 0 0 $X=286810 $Y=211310
X905 2 MASCO__Y15 $T=286810 213310 0 0 $X=286810 $Y=213310
X906 2 MASCO__Y15 $T=286810 215310 0 0 $X=286810 $Y=215310
X907 2 MASCO__Y15 $T=294810 211310 0 0 $X=294810 $Y=211310
X908 2 MASCO__Y15 $T=294810 213310 0 0 $X=294810 $Y=213310
X909 2 MASCO__Y15 $T=294810 215310 0 0 $X=294810 $Y=215310
X910 2 MASCO__Y15 $T=302810 211310 0 0 $X=302810 $Y=211310
X911 2 MASCO__Y15 $T=302810 213310 0 0 $X=302810 $Y=213310
X912 2 MASCO__Y15 $T=302810 215310 0 0 $X=302810 $Y=215310
X913 2 MASCO__Y15 $T=310810 211310 0 0 $X=310810 $Y=211310
X914 2 MASCO__Y15 $T=310810 213310 0 0 $X=310810 $Y=213310
X915 2 MASCO__Y15 $T=310810 215310 0 0 $X=310810 $Y=215310
X916 2 MASCO__Y15 $T=318810 211310 0 0 $X=318810 $Y=211310
X917 2 MASCO__Y15 $T=318810 213310 0 0 $X=318810 $Y=213310
X918 2 MASCO__Y15 $T=318810 215310 0 0 $X=318810 $Y=215310
X919 2 MASCO__Y15 $T=326810 211310 0 0 $X=326810 $Y=211310
X920 2 MASCO__Y15 $T=326810 213310 0 0 $X=326810 $Y=213310
X921 2 MASCO__Y15 $T=326810 215310 0 0 $X=326810 $Y=215310
X922 2 MASCO__Y15 $T=334810 211310 0 0 $X=334810 $Y=211310
X923 2 MASCO__Y15 $T=334810 213310 0 0 $X=334810 $Y=213310
X924 2 MASCO__Y15 $T=334810 215310 0 0 $X=334810 $Y=215310
X925 2 MASCO__Y15 $T=342810 211310 0 0 $X=342810 $Y=211310
X926 2 MASCO__Y15 $T=342810 213310 0 0 $X=342810 $Y=213310
X927 2 MASCO__Y15 $T=342810 215310 0 0 $X=342810 $Y=215310
X928 2 MASCO__Y15 $T=350810 211310 0 0 $X=350810 $Y=211310
X929 2 MASCO__Y15 $T=350810 213310 0 0 $X=350810 $Y=213310
X930 2 MASCO__Y15 $T=350810 215310 0 0 $X=350810 $Y=215310
X931 2 MASCO__Y15 $T=358810 211310 0 0 $X=358810 $Y=211310
X932 2 MASCO__Y15 $T=358810 213310 0 0 $X=358810 $Y=213310
X933 2 MASCO__Y15 $T=358810 215310 0 0 $X=358810 $Y=215310
X934 2 MASCO__Y15 $T=366810 211310 0 0 $X=366810 $Y=211310
X935 2 MASCO__Y15 $T=366810 213310 0 0 $X=366810 $Y=213310
X936 2 MASCO__Y15 $T=366810 215310 0 0 $X=366810 $Y=215310
X937 2 MASCO__Y16 $T=271810 228310 0 0 $X=271810 $Y=228310
X938 2 MASCO__Y16 $T=279810 228310 0 0 $X=279810 $Y=228310
X939 2 MASCO__Y16 $T=287810 228310 0 0 $X=287810 $Y=228310
X940 2 MASCO__Y16 $T=295810 228310 0 0 $X=295810 $Y=228310
X941 2 MASCO__Y16 $T=303810 228310 0 0 $X=303810 $Y=228310
X942 2 MASCO__Y16 $T=311810 228310 0 0 $X=311810 $Y=228310
X943 2 MASCO__Y16 $T=319810 228310 0 0 $X=319810 $Y=228310
X944 2 MASCO__Y16 $T=327810 228310 0 0 $X=327810 $Y=228310
X945 2 MASCO__Y16 $T=335810 228310 0 0 $X=335810 $Y=228310
X946 2 MASCO__Y16 $T=343810 228310 0 0 $X=343810 $Y=228310
X947 2 MASCO__Y16 $T=351810 228310 0 0 $X=351810 $Y=228310
X948 2 MASCO__Y16 $T=359810 228310 0 0 $X=359810 $Y=228310
X949 2 MASCO__Y16 $T=367810 228310 0 0 $X=367810 $Y=228310
X950 9 MASCO__Y16 $T=378495 155110 0 0 $X=378495 $Y=155110
X951 2 MASCO__Y17 $T=270810 217310 0 0 $X=270810 $Y=217310
X952 2 MASCO__Y17 $T=282810 217310 0 0 $X=282810 $Y=217310
X953 2 MASCO__Y17 $T=294810 217310 0 0 $X=294810 $Y=217310
X954 2 MASCO__Y17 $T=306810 217310 0 0 $X=306810 $Y=217310
X955 2 MASCO__Y17 $T=318810 217310 0 0 $X=318810 $Y=217310
X956 2 MASCO__Y17 $T=330810 217310 0 0 $X=330810 $Y=217310
X957 2 MASCO__Y17 $T=342810 217310 0 0 $X=342810 $Y=217310
X958 2 MASCO__Y17 $T=354810 217310 0 0 $X=354810 $Y=217310
X959 2 MASCO__Y18 $T=270810 209070 0 0 $X=270810 $Y=209070
X960 2 MASCO__Y18 $T=276810 209070 0 0 $X=276810 $Y=209070
X961 2 MASCO__Y18 $T=282810 209070 0 0 $X=282810 $Y=209070
X962 2 MASCO__Y18 $T=288810 209070 0 0 $X=288810 $Y=209070
X963 2 MASCO__Y18 $T=294810 209070 0 0 $X=294810 $Y=209070
X964 2 MASCO__Y18 $T=300810 209070 0 0 $X=300810 $Y=209070
X965 2 MASCO__Y18 $T=306810 209070 0 0 $X=306810 $Y=209070
X966 2 MASCO__Y18 $T=312810 209070 0 0 $X=312810 $Y=209070
X967 2 MASCO__Y18 $T=318810 209070 0 0 $X=318810 $Y=209070
X968 2 MASCO__Y18 $T=324810 209070 0 0 $X=324810 $Y=209070
X969 2 MASCO__Y18 $T=330810 209070 0 0 $X=330810 $Y=209070
X970 2 MASCO__Y18 $T=336810 209070 0 0 $X=336810 $Y=209070
X971 2 MASCO__Y18 $T=342810 209070 0 0 $X=342810 $Y=209070
X972 2 MASCO__Y18 $T=348810 209070 0 0 $X=348810 $Y=209070
X973 2 MASCO__Y18 $T=354810 209070 0 0 $X=354810 $Y=209070
X974 2 MASCO__Y18 $T=360810 209070 0 0 $X=360810 $Y=209070
X975 2 MASCO__Y18 $T=366810 209070 0 0 $X=366810 $Y=209070
X976 9 MASCO__Y19 $T=233495 172110 0 0 $X=233495 $Y=172110
X977 9 MASCO__Y19 $T=245495 172110 0 0 $X=245495 $Y=172110
X978 9 MASCO__Y19 $T=269495 172110 0 0 $X=269495 $Y=172110
X979 9 MASCO__Y19 $T=281495 172110 0 0 $X=281495 $Y=172110
X980 9 MASCO__Y19 $T=293495 172110 0 0 $X=293495 $Y=172110
X981 9 MASCO__Y19 $T=305495 172110 0 0 $X=305495 $Y=172110
X982 9 MASCO__Y19 $T=317495 172110 0 0 $X=317495 $Y=172110
X983 9 MASCO__Y19 $T=329495 172110 0 0 $X=329495 $Y=172110
X984 9 MASCO__Y19 $T=341495 172110 0 0 $X=341495 $Y=172110
X985 9 MASCO__Y19 $T=353495 172110 0 0 $X=353495 $Y=172110
D0 1 5 p_dnw AREA=3.39001e-11 PJ=3.421e-05 perimeter=3.421e-05 $X=17815 $Y=113330 $dt=4
D1 1 5 p_dnw3 AREA=2.49e-11 PJ=0 perimeter=0 $X=19030 $Y=114495 $dt=9
.ends MASCO__P3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: hvswitch8                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt hvswitch8 4 8 10 5 3 9 7 6 1
** N=10 EP=9 FDC=433
X0 1 2 3 4 MASCO__H1 $T=0 0 0 0 $X=222710 $Y=91520
X1 1 5 6 3 2 4 MASCO__P2 $T=0 0 0 0 $X=5800 $Y=7480
X2 1 6 2 5 7 8 9 10 3 4 MASCO__P3 $T=0 0 0 0 $X=5800 $Y=102950
.ends hvswitch8
